// Generated from iroha-0.0.1.

// SRAM(2 port(s))
module SRAM_4_32_2(clk, rst, addr_0_i, rdata_0_o, wdata_0_i, write_en_0_i, addr_1_i, rdata_1_o, wdata_1_i, write_en_1_i);
  input clk;
  input rst;
  input [3:0] addr_0_i;
  output [31:0] rdata_0_o;
  input [31:0] wdata_0_i;
  input write_en_0_i;

  reg [31:0] rdata_0_o;

  input [3:0] addr_1_i;
  output [31:0] rdata_1_o;
  input [31:0] wdata_1_i;
  input write_en_1_i;

  reg [31:0] rdata_1_o;

  reg [31:0] data [0:15];

  always @(posedge clk) begin
    if (rst) begin
    end else begin
      if (write_en_0_i) begin
        data[addr_0_i] <= wdata_0_i;
      end
      if (write_en_1_i) begin
        data[addr_1_i] <= wdata_1_i;
      end
    end
  end
  // Read
  always @(addr_0_i or clk) begin
    rdata_0_o = data[addr_0_i];
  end
  always @(addr_1_i or clk) begin
    rdata_1_o = data[addr_1_i];
  end
endmodule


// SRAM(1 port(s))
module SRAM_3_32(clk, rst, addr_i, rdata_o, wdata_i, write_en_i);
  input clk;
  input rst;
  input [2:0] addr_i;
  output [31:0] rdata_o;
  input [31:0] wdata_i;
  input write_en_i;

  reg [31:0] rdata_o;

  reg [31:0] data [0:7];

  always @(posedge clk) begin
    if (rst) begin
      data[0] <= 0;
      data[1] <= 0;
      data[2] <= 0;
      data[3] <= 0;
      data[4] <= 0;
      data[5] <= 0;
      data[6] <= 0;
      data[7] <= 0;
    end else begin
      if (write_en_i) begin
        data[addr_i] <= wdata_i;
      end
    end
  end
  // Read
  always @(addr_i or clk) begin
    rdata_o = data[addr_i];
  end
endmodule


// SRAM(1 port(s))
module SRAM_6_32(clk, rst, addr_i, rdata_o, wdata_i, write_en_i);
  input clk;
  input rst;
  input [5:0] addr_i;
  output [31:0] rdata_o;
  input [31:0] wdata_i;
  input write_en_i;

  reg [31:0] rdata_o;

  reg [31:0] data [0:63];

  always @(posedge clk) begin
    if (rst) begin
      data[0] <= 1116352408;
      data[1] <= 1899447441;
      data[2] <= 3049323471;
      data[3] <= 3921009573;
      data[4] <= 961987163;
      data[5] <= 1508970993;
      data[6] <= 2453635748;
      data[7] <= 2870763221;
      data[8] <= 3624381080;
      data[9] <= 310598401;
      data[10] <= 607225278;
      data[11] <= 1426881987;
      data[12] <= 1925078388;
      data[13] <= 2162078206;
      data[14] <= 2614888103;
      data[15] <= 3248222580;
      data[16] <= 3835390401;
      data[17] <= 4022224774;
      data[18] <= 264347078;
      data[19] <= 604807628;
      data[20] <= 770255983;
      data[21] <= 1249150122;
      data[22] <= 1555081692;
      data[23] <= 1996064986;
      data[24] <= 2554220882;
      data[25] <= 2821834349;
      data[26] <= 2952996808;
      data[27] <= 3210313671;
      data[28] <= 3336571891;
      data[29] <= 3584528711;
      data[30] <= 113926993;
      data[31] <= 338241895;
      data[32] <= 666307205;
      data[33] <= 773529912;
      data[34] <= 1294757372;
      data[35] <= 1396182291;
      data[36] <= 1695183700;
      data[37] <= 1986661051;
      data[38] <= 2177026350;
      data[39] <= 2456956037;
      data[40] <= 2730485921;
      data[41] <= 2820302411;
      data[42] <= 3259730800;
      data[43] <= 3345764771;
      data[44] <= 3516065817;
      data[45] <= 3600352804;
      data[46] <= 4094571909;
      data[47] <= 275423344;
      data[48] <= 430227734;
      data[49] <= 506948616;
      data[50] <= 659060556;
      data[51] <= 883997877;
      data[52] <= 958139571;
      data[53] <= 1322822218;
      data[54] <= 1537002063;
      data[55] <= 1747873779;
      data[56] <= 1955562222;
      data[57] <= 2024104815;
      data[58] <= 2227730452;
      data[59] <= 2361852424;
      data[60] <= 2428436474;
      data[61] <= 2756734187;
      data[62] <= 3204031479;
      data[63] <= 3329325298;
    end else begin
      if (write_en_i) begin
        data[addr_i] <= wdata_i;
      end
    end
  end
  // Read
  always @(addr_i or clk) begin
    rdata_o = data[addr_i];
  end
endmodule

module axi_master_controller_a4rd32(clk, rst, sram_addr, sram_wdata, sram_wen, sram_rdata, sram_EXCLUSIVE, sram_req, sram_ack, addr, len, start, wen, req, ack, ARADDR, ARVALID, ARREADY, ARLEN, ARSIZE, RVALID, RDATA, RREADY, RLAST, AWADDR, AWVALID, AWREADY, AWLEN, AWSIZE, WVALID, WREADY, WDATA, WLAST, BVALID, BREADY, BRESP);
  input clk;
  input rst;
  output [3:0] sram_addr;
  output [31:0] sram_wdata;
  output sram_wen;
  input [31:0] sram_rdata;
  input sram_EXCLUSIVE;
  output sram_req;
  input sram_ack;
  input [31:0] addr;
  input [3:0] len;
  input [3:0] start;
  input wen;
  input req;
  output ack;
  output [31:0] ARADDR;
  output ARVALID;
  input ARREADY;
  output [7:0] ARLEN;
  output [2:0] ARSIZE;
  input RVALID;
  input [31:0] RDATA;
  output RREADY;
  input RLAST;
  output [31:0] AWADDR;
  output AWVALID;
  input AWREADY;
  output [7:0] AWLEN;
  output [2:0] AWSIZE;
  output WVALID;
  input WREADY;
  output [31:0] WDATA;
  output WLAST;
  input BVALID;
  output BREADY;
  input [1:0] BRESP;
  reg [3:0] sram_addr;
  reg [31:0] sram_wdata;
  reg sram_wen;
  reg sram_req;
  reg ack;
  reg [31:0] ARADDR;
  reg ARVALID;
  reg [7:0] ARLEN;
  reg [2:0] ARSIZE;
  reg RREADY;
  reg [31:0] AWADDR;
  reg AWVALID;
  reg [7:0] AWLEN;
  reg [2:0] AWSIZE;
  reg WVALID;
  reg [31:0] WDATA;
  reg WLAST;
  reg BREADY;

  `define S_IDLE 0
  `define S_ADDR_WAIT 1
  `define S_READ_DATA 2
  `define S_READ_DATA_WAIT 3
  reg [2:0] st;

  reg [4:0] ridx;
  reg read_last;

  always @(posedge clk) begin
    if (rst) begin
      ack <= 0;
      sram_req <= 0;
      sram_wen <= 0;
      st <= `S_IDLE;
      ARADDR <= 0;
      ARVALID <= 0;
      ARLEN <= 0;
      ARSIZE <= 0;
      RREADY <= 0;
      AWADDR <= 0;
      AWVALID <= 0;
      AWLEN <= 0;
      AWSIZE <= 0;
      WVALID <= 0;
      WDATA <= 0;
      WLAST <= 0;
      BREADY <= 0;
    end else begin
      if (sram_EXCLUSIVE) begin
        sram_wen <= (st == `S_READ_DATA && RVALID);
      end
      case (st)
        `S_IDLE: begin
          ack <= 0;
          if (req && !ack) begin
            ridx <= 0;
            st <= `S_ADDR_WAIT;
            ARVALID <= 1;
            ARADDR <= addr;
            ARLEN <= len;
            ARSIZE <= 2;
          end
        end
        `S_ADDR_WAIT: begin
          ack <= 0;
          if (ARREADY) begin
            st <= `S_READ_DATA;
            ARVALID <= 0;
            RREADY <= 1;
          end
        end
        `S_READ_DATA: begin
          if (RVALID) begin
            sram_addr <= start + ridx;
            sram_wdata <= RDATA;
            ridx <= ridx + 1;
            if (sram_EXCLUSIVE) begin
              if (RLAST) begin
                RREADY <= 0;
                ack <= 1;
                st <= `S_IDLE;
              end
            end else begin
              st <= `S_READ_DATA_WAIT;
              sram_req <= 1;
              sram_wen <= 1;
              RREADY <= 0;
              read_last <= RLAST;
            end
          end
        end
        `S_READ_DATA_WAIT: begin
          if (sram_ack) begin
            sram_req <= 0;
            sram_wen <= 0;
            if (read_last) begin
              ack <= 1;
              st <= `S_IDLE;
            end else begin
              st <= `S_READ_DATA;
              RREADY <= 1;
            end
          end
        end
      endcase
    end
  end
endmodule

// Module 1;
module main(clk, rst, buf_ARADDR, buf_ARVALID, buf_ARREADY, buf_ARLEN, buf_ARSIZE, buf_RVALID, buf_RDATA, buf_RREADY, buf_RLAST, buf_AWADDR, buf_AWVALID, buf_AWREADY, buf_AWLEN, buf_AWSIZE, buf_WVALID, buf_WREADY, buf_WDATA, buf_WLAST, buf_BVALID, buf_BREADY, buf_BRESP, sha256_req_valid, sha256_req_ready, sha256_req_busy, sha256_res_valid, sha256_res_ready, sha256_req_0, sha256_req_1, sha256_res_0);
  input clk;
  input rst;
  output [31:0] buf_ARADDR;
  output buf_ARVALID;
  input buf_ARREADY;
  output [7:0] buf_ARLEN;
  output [2:0] buf_ARSIZE;
  input buf_RVALID;
  input [31:0] buf_RDATA;
  output buf_RREADY;
  input buf_RLAST;
  output [31:0] buf_AWADDR;
  output buf_AWVALID;
  input buf_AWREADY;
  output [7:0] buf_AWLEN;
  output [2:0] buf_AWSIZE;
  output buf_WVALID;
  input buf_WREADY;
  output [31:0] buf_WDATA;
  output buf_WLAST;
  input buf_BVALID;
  output buf_BREADY;
  input [1:0] buf_BRESP;
  input sha256_req_valid;
  output sha256_req_ready;
  output sha256_req_busy;
  output sha256_res_valid;
  input sha256_res_ready;
  input [31:0] sha256_req_0;
  input [31:0] sha256_req_1;
  output [255:0] sha256_res_0;
  reg sha256_req_ready;
  reg sha256_req_busy;
  reg sha256_res_valid;
  reg [255:0] sha256_res_0;

  // State decls
  // state names
  `define S_1_1 1
  `define S_1_2 2
  reg [1:0] st_1;

  // state names
  `define S_2_1 1
  `define S_2_6 6
  `define S_2_7 7
  `define S_2_8 8
  `define S_2_9 9
  `define S_2_13 13
  `define S_2_19 19
  `define S_2_20 20
  `define S_2_21 21
  `define S_2_23 23
  `define S_2_26 26
  `define S_2_2 2
  `define S_2_30 30
  `define S_2_3 3
  `define S_2_31 31
  `define S_2_35 35
  `define S_2_4 4
  `define S_2_36 36
  `define S_2_40 40
  `define S_2_5 5
  `define S_2_41 41
  `define S_2_45 45
  `define S_2_10 10
  `define S_2_46 46
  `define S_2_50 50
  `define S_2_11 11
  `define S_2_51 51
  `define S_2_55 55
  `define S_2_12 12
  `define S_2_56 56
  `define S_2_60 60
  `define S_2_14 14
  `define S_2_61 61
  `define S_2_62 62
  `define S_2_66 66
  `define S_2_72 72
  `define S_2_77 77
  `define S_2_82 82
  `define S_2_87 87
  `define S_2_92 92
  `define S_2_97 97
  `define S_2_102 102
  `define S_2_107 107
  `define S_2_113 113
  `define S_2_114 114
  `define S_2_115 115
  `define S_2_116 116
  `define S_2_117 117
  `define S_2_120 120
  `define S_2_121 121
  `define S_2_122 122
  `define S_2_125 125
  `define S_2_126 126
  `define S_2_128 128
  `define S_2_129 129
  `define S_2_130 130
  `define S_2_131 131
  `define S_2_132 132
  `define S_2_133 133
  `define S_2_135 135
  `define S_2_138 138
  `define S_2_15 15
  `define S_2_139 139
  `define S_2_140 140
  `define S_2_142 142
  `define S_2_145 145
  `define S_2_16 16
  `define S_2_146 146
  `define S_2_149 149
  `define S_2_152 152
  `define S_2_17 17
  `define S_2_153 153
  `define S_2_154 154
  `define S_2_155 155
  `define S_2_157 157
  `define S_2_160 160
  `define S_2_18 18
  `define S_2_161 161
  `define S_2_164 164
  `define S_2_165 165
  `define S_2_167 167
  `define S_2_170 170
  `define S_2_22 22
  `define S_2_171 171
  `define S_2_175 175
  `define S_2_24 24
  `define S_2_176 176
  `define S_2_180 180
  `define S_2_25 25
  `define S_2_181 181
  `define S_2_185 185
  `define S_2_27 27
  `define S_2_186 186
  `define S_2_190 190
  `define S_2_28 28
  `define S_2_191 191
  `define S_2_195 195
  `define S_2_29 29
  `define S_2_196 196
  `define S_2_200 200
  `define S_2_32 32
  `define S_2_201 201
  `define S_2_205 205
  `define S_2_33 33
  `define S_2_206 206
  `define S_2_208 208
  `define S_2_209 209
  `define S_2_210 210
  `define S_2_211 211
  `define S_2_212 212
  `define S_2_213 213
  `define S_2_214 214
  `define S_2_216 216
  `define S_2_217 217
  `define S_2_219 219
  `define S_2_222 222
  `define S_2_34 34
  `define S_2_223 223
  `define S_2_227 227
  `define S_2_231 231
  `define S_2_37 37
  `define S_2_232 232
  `define S_2_236 236
  `define S_2_240 240
  `define S_2_38 38
  `define S_2_241 241
  `define S_2_245 245
  `define S_2_249 249
  `define S_2_39 39
  `define S_2_250 250
  `define S_2_254 254
  `define S_2_258 258
  `define S_2_42 42
  `define S_2_259 259
  `define S_2_263 263
  `define S_2_267 267
  `define S_2_43 43
  `define S_2_268 268
  `define S_2_272 272
  `define S_2_276 276
  `define S_2_44 44
  `define S_2_277 277
  `define S_2_281 281
  `define S_2_285 285
  `define S_2_47 47
  `define S_2_286 286
  `define S_2_290 290
  `define S_2_297 297
  `define S_2_300 300
  `define S_2_301 301
  `define S_2_304 304
  `define S_2_305 305
  `define S_2_308 308
  `define S_2_309 309
  `define S_2_310 310
  `define S_2_317 317
  `define S_2_318 318
  `define S_2_320 320
  `define S_2_321 321
  `define S_2_322 322
  `define S_2_324 324
  `define S_2_325 325
  `define S_2_326 326
  `define S_2_334 334
  `define S_2_337 337
  `define S_2_338 338
  `define S_2_339 339
  `define S_2_347 347
  `define S_2_350 350
  `define S_2_351 351
  `define S_2_352 352
  `define S_2_359 359
  `define S_2_360 360
  `define S_2_362 362
  `define S_2_363 363
  `define S_2_364 364
  `define S_2_366 366
  `define S_2_367 367
  `define S_2_368 368
  `define S_2_376 376
  `define S_2_379 379
  `define S_2_380 380
  `define S_2_381 381
  `define S_2_389 389
  `define S_2_392 392
  `define S_2_393 393
  `define S_2_394 394
  `define S_2_401 401
  `define S_2_402 402
  `define S_2_403 403
  `define S_2_405 405
  `define S_2_406 406
  `define S_2_407 407
  `define S_2_410 410
  `define S_2_48 48
  `define S_2_411 411
  `define S_2_414 414
  `define S_2_49 49
  `define S_2_415 415
  `define S_2_416 416
  `define S_2_418 418
  `define S_2_419 419
  `define S_2_421 421
  `define S_2_422 422
  `define S_2_423 423
  `define S_2_424 424
  `define S_2_425 425
  `define S_2_426 426
  `define S_2_427 427
  `define S_2_428 428
  `define S_2_430 430
  `define S_2_431 431
  `define S_2_432 432
  `define S_2_434 434
  `define S_2_435 435
  `define S_2_436 436
  `define S_2_438 438
  `define S_2_441 441
  `define S_2_52 52
  `define S_2_442 442
  `define S_2_444 444
  `define S_2_447 447
  `define S_2_53 53
  `define S_2_448 448
  `define S_2_449 449
  `define S_2_451 451
  `define S_2_452 452
  `define S_2_454 454
  `define S_2_455 455
  `define S_2_456 456
  `define S_2_457 457
  `define S_2_458 458
  `define S_2_459 459
  `define S_2_460 460
  `define S_2_461 461
  `define S_2_463 463
  `define S_2_464 464
  `define S_2_465 465
  `define S_2_467 467
  `define S_2_468 468
  `define S_2_469 469
  `define S_2_471 471
  `define S_2_474 474
  `define S_2_54 54
  `define S_2_475 475
  `define S_2_477 477
  `define S_2_480 480
  `define S_2_57 57
  `define S_2_481 481
  `define S_2_482 482
  `define S_2_484 484
  `define S_2_485 485
  `define S_2_487 487
  `define S_2_488 488
  `define S_2_489 489
  `define S_2_490 490
  `define S_2_491 491
  `define S_2_492 492
  `define S_2_493 493
  `define S_2_494 494
  `define S_2_496 496
  `define S_2_497 497
  `define S_2_498 498
  `define S_2_500 500
  `define S_2_501 501
  `define S_2_502 502
  `define S_2_504 504
  `define S_2_507 507
  `define S_2_58 58
  `define S_2_508 508
  `define S_2_510 510
  `define S_2_513 513
  `define S_2_59 59
  `define S_2_514 514
  `define S_2_515 515
  `define S_2_517 517
  `define S_2_518 518
  `define S_2_520 520
  `define S_2_521 521
  `define S_2_522 522
  `define S_2_523 523
  `define S_2_524 524
  `define S_2_525 525
  `define S_2_526 526
  `define S_2_527 527
  `define S_2_529 529
  `define S_2_530 530
  `define S_2_531 531
  `define S_2_533 533
  `define S_2_534 534
  `define S_2_535 535
  `define S_2_537 537
  `define S_2_540 540
  `define S_2_63 63
  `define S_2_541 541
  `define S_2_543 543
  `define S_2_546 546
  `define S_2_64 64
  `define S_2_547 547
  `define S_2_548 548
  `define S_2_550 550
  `define S_2_551 551
  `define S_2_553 553
  `define S_2_554 554
  `define S_2_555 555
  `define S_2_556 556
  `define S_2_557 557
  `define S_2_558 558
  `define S_2_559 559
  `define S_2_560 560
  `define S_2_562 562
  `define S_2_563 563
  `define S_2_564 564
  `define S_2_566 566
  `define S_2_567 567
  `define S_2_568 568
  `define S_2_570 570
  `define S_2_573 573
  `define S_2_65 65
  `define S_2_574 574
  `define S_2_576 576
  `define S_2_579 579
  `define S_2_67 67
  `define S_2_580 580
  `define S_2_581 581
  `define S_2_583 583
  `define S_2_584 584
  `define S_2_586 586
  `define S_2_587 587
  `define S_2_588 588
  `define S_2_589 589
  `define S_2_590 590
  `define S_2_591 591
  `define S_2_592 592
  `define S_2_593 593
  `define S_2_595 595
  `define S_2_596 596
  `define S_2_597 597
  `define S_2_599 599
  `define S_2_600 600
  `define S_2_601 601
  `define S_2_603 603
  `define S_2_606 606
  `define S_2_68 68
  `define S_2_607 607
  `define S_2_609 609
  `define S_2_612 612
  `define S_2_69 69
  `define S_2_613 613
  `define S_2_614 614
  `define S_2_616 616
  `define S_2_617 617
  `define S_2_619 619
  `define S_2_620 620
  `define S_2_621 621
  `define S_2_622 622
  `define S_2_623 623
  `define S_2_624 624
  `define S_2_625 625
  `define S_2_626 626
  `define S_2_628 628
  `define S_2_629 629
  `define S_2_630 630
  `define S_2_632 632
  `define S_2_633 633
  `define S_2_634 634
  `define S_2_636 636
  `define S_2_639 639
  `define S_2_70 70
  `define S_2_640 640
  `define S_2_642 642
  `define S_2_645 645
  `define S_2_71 71
  `define S_2_646 646
  `define S_2_647 647
  `define S_2_649 649
  `define S_2_650 650
  `define S_2_652 652
  `define S_2_653 653
  `define S_2_654 654
  `define S_2_655 655
  `define S_2_656 656
  `define S_2_657 657
  `define S_2_658 658
  `define S_2_659 659
  `define S_2_660 660
  `define S_2_661 661
  `define S_2_662 662
  `define S_2_663 663
  `define S_2_664 664
  `define S_2_665 665
  `define S_2_666 666
  `define S_2_667 667
  `define S_2_674 674
  `define S_2_675 675
  `define S_2_677 677
  `define S_2_678 678
  `define S_2_679 679
  `define S_2_681 681
  `define S_2_682 682
  `define S_2_683 683
  `define S_2_684 684
  `define S_2_692 692
  `define S_2_695 695
  `define S_2_696 696
  `define S_2_697 697
  `define S_2_705 705
  `define S_2_708 708
  `define S_2_709 709
  `define S_2_710 710
  `define S_2_718 718
  `define S_2_721 721
  `define S_2_722 722
  `define S_2_723 723
  `define S_2_729 729
  `define S_2_730 730
  `define S_2_731 731
  `define S_2_732 732
  `define S_2_739 739
  `define S_2_740 740
  `define S_2_742 742
  `define S_2_743 743
  `define S_2_744 744
  `define S_2_746 746
  `define S_2_747 747
  `define S_2_748 748
  `define S_2_749 749
  `define S_2_757 757
  `define S_2_760 760
  `define S_2_761 761
  `define S_2_762 762
  `define S_2_770 770
  `define S_2_773 773
  `define S_2_774 774
  `define S_2_775 775
  `define S_2_783 783
  `define S_2_786 786
  `define S_2_787 787
  `define S_2_788 788
  `define S_2_794 794
  `define S_2_795 795
  `define S_2_796 796
  `define S_2_797 797
  `define S_2_798 798
  `define S_2_805 805
  `define S_2_806 806
  `define S_2_808 808
  `define S_2_809 809
  `define S_2_810 810
  `define S_2_812 812
  `define S_2_813 813
  `define S_2_814 814
  `define S_2_815 815
  `define S_2_823 823
  `define S_2_826 826
  `define S_2_827 827
  `define S_2_828 828
  `define S_2_836 836
  `define S_2_839 839
  `define S_2_840 840
  `define S_2_841 841
  `define S_2_849 849
  `define S_2_852 852
  `define S_2_853 853
  `define S_2_854 854
  `define S_2_860 860
  `define S_2_861 861
  `define S_2_862 862
  `define S_2_863 863
  `define S_2_870 870
  `define S_2_871 871
  `define S_2_873 873
  `define S_2_874 874
  `define S_2_875 875
  `define S_2_877 877
  `define S_2_878 878
  `define S_2_879 879
  `define S_2_880 880
  `define S_2_888 888
  `define S_2_891 891
  `define S_2_892 892
  `define S_2_893 893
  `define S_2_901 901
  `define S_2_904 904
  `define S_2_905 905
  `define S_2_906 906
  `define S_2_914 914
  `define S_2_917 917
  `define S_2_918 918
  `define S_2_919 919
  `define S_2_925 925
  `define S_2_926 926
  `define S_2_927 927
  `define S_2_928 928
  `define S_2_929 929
  `define S_2_936 936
  `define S_2_937 937
  `define S_2_939 939
  `define S_2_940 940
  `define S_2_941 941
  `define S_2_943 943
  `define S_2_944 944
  `define S_2_945 945
  `define S_2_946 946
  `define S_2_954 954
  `define S_2_957 957
  `define S_2_958 958
  `define S_2_959 959
  `define S_2_967 967
  `define S_2_970 970
  `define S_2_971 971
  `define S_2_972 972
  `define S_2_980 980
  `define S_2_983 983
  `define S_2_984 984
  `define S_2_985 985
  `define S_2_991 991
  `define S_2_992 992
  `define S_2_993 993
  `define S_2_994 994
  `define S_2_1001 1001
  `define S_2_1002 1002
  `define S_2_1004 1004
  `define S_2_1005 1005
  `define S_2_1006 1006
  `define S_2_1008 1008
  `define S_2_1009 1009
  `define S_2_1010 1010
  `define S_2_1011 1011
  `define S_2_1019 1019
  `define S_2_1022 1022
  `define S_2_1023 1023
  `define S_2_1024 1024
  `define S_2_1032 1032
  `define S_2_1035 1035
  `define S_2_1036 1036
  `define S_2_1037 1037
  `define S_2_1045 1045
  `define S_2_1048 1048
  `define S_2_1049 1049
  `define S_2_1050 1050
  `define S_2_1056 1056
  `define S_2_1057 1057
  `define S_2_1058 1058
  `define S_2_1059 1059
  `define S_2_1060 1060
  `define S_2_1067 1067
  `define S_2_1068 1068
  `define S_2_1070 1070
  `define S_2_1071 1071
  `define S_2_1072 1072
  `define S_2_1074 1074
  `define S_2_1075 1075
  `define S_2_1076 1076
  `define S_2_1077 1077
  `define S_2_1085 1085
  `define S_2_1088 1088
  `define S_2_1089 1089
  `define S_2_1090 1090
  `define S_2_1098 1098
  `define S_2_1101 1101
  `define S_2_1102 1102
  `define S_2_1103 1103
  `define S_2_1111 1111
  `define S_2_1114 1114
  `define S_2_1115 1115
  `define S_2_1116 1116
  `define S_2_1122 1122
  `define S_2_1123 1123
  `define S_2_1124 1124
  `define S_2_1125 1125
  `define S_2_1132 1132
  `define S_2_1133 1133
  `define S_2_1135 1135
  `define S_2_1136 1136
  `define S_2_1137 1137
  `define S_2_1139 1139
  `define S_2_1140 1140
  `define S_2_1141 1141
  `define S_2_1142 1142
  `define S_2_1150 1150
  `define S_2_1153 1153
  `define S_2_1154 1154
  `define S_2_1155 1155
  `define S_2_1163 1163
  `define S_2_1166 1166
  `define S_2_1167 1167
  `define S_2_1168 1168
  `define S_2_1176 1176
  `define S_2_1179 1179
  `define S_2_1180 1180
  `define S_2_1181 1181
  `define S_2_1187 1187
  `define S_2_1188 1188
  `define S_2_1189 1189
  `define S_2_1190 1190
  `define S_2_1191 1191
  `define S_2_1198 1198
  `define S_2_1199 1199
  `define S_2_1201 1201
  `define S_2_1202 1202
  `define S_2_1203 1203
  `define S_2_1205 1205
  `define S_2_1206 1206
  `define S_2_1207 1207
  `define S_2_1208 1208
  `define S_2_1216 1216
  `define S_2_1219 1219
  `define S_2_1220 1220
  `define S_2_1221 1221
  `define S_2_1229 1229
  `define S_2_1232 1232
  `define S_2_1233 1233
  `define S_2_1234 1234
  `define S_2_1242 1242
  `define S_2_1245 1245
  `define S_2_1246 1246
  `define S_2_1247 1247
  `define S_2_1253 1253
  `define S_2_1254 1254
  `define S_2_1255 1255
  `define S_2_1256 1256
  `define S_2_1263 1263
  `define S_2_1264 1264
  `define S_2_1266 1266
  `define S_2_1267 1267
  `define S_2_1268 1268
  `define S_2_1270 1270
  `define S_2_1271 1271
  `define S_2_1272 1272
  `define S_2_1273 1273
  `define S_2_1281 1281
  `define S_2_1284 1284
  `define S_2_1285 1285
  `define S_2_1286 1286
  `define S_2_1294 1294
  `define S_2_1297 1297
  `define S_2_1298 1298
  `define S_2_1299 1299
  `define S_2_1307 1307
  `define S_2_1310 1310
  `define S_2_1311 1311
  `define S_2_1312 1312
  `define S_2_1318 1318
  `define S_2_1319 1319
  `define S_2_1320 1320
  `define S_2_1321 1321
  `define S_2_1322 1322
  `define S_2_1329 1329
  `define S_2_1330 1330
  `define S_2_1332 1332
  `define S_2_1333 1333
  `define S_2_1334 1334
  `define S_2_1336 1336
  `define S_2_1337 1337
  `define S_2_1338 1338
  `define S_2_1339 1339
  `define S_2_1347 1347
  `define S_2_1350 1350
  `define S_2_1351 1351
  `define S_2_1352 1352
  `define S_2_1360 1360
  `define S_2_1363 1363
  `define S_2_1364 1364
  `define S_2_1365 1365
  `define S_2_1373 1373
  `define S_2_1376 1376
  `define S_2_1377 1377
  `define S_2_1378 1378
  `define S_2_1384 1384
  `define S_2_1385 1385
  `define S_2_1386 1386
  `define S_2_1387 1387
  `define S_2_1394 1394
  `define S_2_1395 1395
  `define S_2_1397 1397
  `define S_2_1398 1398
  `define S_2_1399 1399
  `define S_2_1401 1401
  `define S_2_1402 1402
  `define S_2_1403 1403
  `define S_2_1404 1404
  `define S_2_1412 1412
  `define S_2_1415 1415
  `define S_2_1416 1416
  `define S_2_1417 1417
  `define S_2_1425 1425
  `define S_2_1428 1428
  `define S_2_1429 1429
  `define S_2_1430 1430
  `define S_2_1438 1438
  `define S_2_1441 1441
  `define S_2_1442 1442
  `define S_2_1443 1443
  `define S_2_1449 1449
  `define S_2_1450 1450
  `define S_2_1451 1451
  `define S_2_1452 1452
  `define S_2_1453 1453
  `define S_2_1460 1460
  `define S_2_1461 1461
  `define S_2_1463 1463
  `define S_2_1464 1464
  `define S_2_1465 1465
  `define S_2_1467 1467
  `define S_2_1468 1468
  `define S_2_1469 1469
  `define S_2_1470 1470
  `define S_2_1478 1478
  `define S_2_1481 1481
  `define S_2_1482 1482
  `define S_2_1483 1483
  `define S_2_1491 1491
  `define S_2_1494 1494
  `define S_2_1495 1495
  `define S_2_1496 1496
  `define S_2_1504 1504
  `define S_2_1507 1507
  `define S_2_1508 1508
  `define S_2_1509 1509
  `define S_2_1515 1515
  `define S_2_1516 1516
  `define S_2_1517 1517
  `define S_2_1518 1518
  `define S_2_1525 1525
  `define S_2_1526 1526
  `define S_2_1528 1528
  `define S_2_1529 1529
  `define S_2_1530 1530
  `define S_2_1532 1532
  `define S_2_1533 1533
  `define S_2_1534 1534
  `define S_2_1535 1535
  `define S_2_1543 1543
  `define S_2_1546 1546
  `define S_2_1547 1547
  `define S_2_1548 1548
  `define S_2_1556 1556
  `define S_2_1559 1559
  `define S_2_1560 1560
  `define S_2_1561 1561
  `define S_2_1569 1569
  `define S_2_1572 1572
  `define S_2_1573 1573
  `define S_2_1574 1574
  `define S_2_1580 1580
  `define S_2_1581 1581
  `define S_2_1582 1582
  `define S_2_1583 1583
  `define S_2_1584 1584
  `define S_2_1591 1591
  `define S_2_1592 1592
  `define S_2_1594 1594
  `define S_2_1595 1595
  `define S_2_1596 1596
  `define S_2_1598 1598
  `define S_2_1599 1599
  `define S_2_1600 1600
  `define S_2_1601 1601
  `define S_2_1609 1609
  `define S_2_1612 1612
  `define S_2_1613 1613
  `define S_2_1614 1614
  `define S_2_1622 1622
  `define S_2_1625 1625
  `define S_2_1626 1626
  `define S_2_1627 1627
  `define S_2_1635 1635
  `define S_2_1638 1638
  `define S_2_1639 1639
  `define S_2_1640 1640
  `define S_2_1646 1646
  `define S_2_1647 1647
  `define S_2_1648 1648
  `define S_2_1649 1649
  `define S_2_1656 1656
  `define S_2_1657 1657
  `define S_2_1659 1659
  `define S_2_1660 1660
  `define S_2_1661 1661
  `define S_2_1663 1663
  `define S_2_1664 1664
  `define S_2_1665 1665
  `define S_2_1666 1666
  `define S_2_1674 1674
  `define S_2_1677 1677
  `define S_2_1678 1678
  `define S_2_1679 1679
  `define S_2_1687 1687
  `define S_2_1690 1690
  `define S_2_1691 1691
  `define S_2_1692 1692
  `define S_2_1700 1700
  `define S_2_1703 1703
  `define S_2_1704 1704
  `define S_2_1705 1705
  `define S_2_1711 1711
  `define S_2_1712 1712
  `define S_2_1713 1713
  `define S_2_1714 1714
  `define S_2_1715 1715
  `define S_2_task_idle 1716
  reg [11:0] st_2;

  // State vars
  // Registers
  reg  [31:0] r__38_335;
  reg  [31:0] arg_15_389;
  reg  [31:0] r1_bswap_16_397;
  reg  [7:0] r5_bswap_17_390;
  reg  [7:0] r8_bswap_18_391;
  reg  [15:0] r4_bswap_19_392;
  reg  [7:0] r11_bswap_20_393;
  reg  [23:0] r3_bswap_21_394;
  reg  [7:0] r14_bswap_22_395;
  reg  [31:0] r2_bswap_23_396;
  reg  [14:0] r6_ror32_17_189_407;
  reg  [31:0] r2_ror32_17_190_408;
  reg  [31:0] arg_186_405;
  reg  [31:0] r1_ror32_17_187_409;
  reg  [16:0] r3_ror32_17_188_406;
  reg  [31:0] arg_196_410;
  reg  [31:0] r1_ror32_19_197_414;
  reg  [18:0] r3_ror32_19_198_411;
  reg  [12:0] r6_ror32_19_199_412;
  reg  [31:0] r2_ror32_19_200_413;
  reg  [31:0] x_233_398;
  reg  [31:0] r1_s1_234_404;
  reg  [31:0] r4_s1_235_399;
  reg  [31:0] r6_s1_236_400;
  reg  [31:0] r3_s1_237_401;
  reg  [31:0] r8_s1_238_402;
  reg  [31:0] r2_s1_239_403;
  reg  [6:0] r3_ror32_7_223_423;
  reg  [24:0] r6_ror32_7_224_424;
  reg  [31:0] arg_221_422;
  reg  [31:0] r1_ror32_7_222_426;
  reg  [31:0] r2_ror32_7_225_425;
  reg  [31:0] arg_191_427;
  reg  [31:0] r1_ror32_18_192_431;
  reg  [17:0] r3_ror32_18_193_428;
  reg  [13:0] r6_ror32_18_194_429;
  reg  [31:0] r2_ror32_18_195_430;
  reg  [31:0] x_226_415;
  reg  [31:0] r1_s0_227_421;
  reg  [31:0] r4_s0_228_416;
  reg  [31:0] r6_s0_229_417;
  reg  [31:0] r3_s0_230_418;
  reg  [31:0] r8_s0_231_419;
  reg  [31:0] r2_s0_232_420;
  reg  [31:0] arg_216_576;
  reg  [31:0] r1_ror32_6_217_580;
  reg  [5:0] r3_ror32_6_218_577;
  reg  [25:0] r6_ror32_6_219_578;
  reg  [31:0] r2_ror32_6_220_579;
  reg  [31:0] arg_176_581;
  reg  [31:0] r1_ror32_11_177_585;
  reg  [10:0] r3_ror32_11_178_582;
  reg  [20:0] r6_ror32_11_179_583;
  reg  [31:0] r2_ror32_11_180_584;
  reg  [31:0] arg_211_586;
  reg  [31:0] r1_ror32_25_212_590;
  reg  [24:0] r3_ror32_25_213_587;
  reg  [6:0] r6_ror32_25_214_588;
  reg  [31:0] r2_ror32_25_215_589;
  reg  [31:0] x_31_569;
  reg  [31:0] r1_e1_32_575;
  reg  [31:0] r4_e1_33_570;
  reg  [31:0] r6_e1_34_571;
  reg  [31:0] r3_e1_35_572;
  reg  [31:0] r8_e1_36_573;
  reg  [31:0] r2_e1_37_574;
  reg  [31:0] x_0_594;
  reg  [31:0] y_1_591;
  reg  [31:0] z_2_592;
  reg  [31:0] r3_Ch_3_597;
  reg  [31:0] r6_Ch_4_593;
  reg  [31:0] r5_Ch_5_595;
  reg  [31:0] r4_Ch_6_596;
  reg  [31:0] arg_201_605;
  reg  [31:0] r1_ror32_2_202_609;
  reg  [1:0] r3_ror32_2_203_606;
  reg  [29:0] r6_ror32_2_204_607;
  reg  [31:0] r2_ror32_2_205_608;
  reg  [31:0] arg_181_610;
  reg  [31:0] r1_ror32_13_182_614;
  reg  [12:0] r3_ror32_13_183_611;
  reg  [18:0] r6_ror32_13_184_612;
  reg  [31:0] r2_ror32_13_185_613;
  reg  [31:0] arg_206_615;
  reg  [31:0] r1_ror32_22_207_619;
  reg  [21:0] r3_ror32_22_208_616;
  reg  [9:0] r6_ror32_22_209_617;
  reg  [31:0] r2_ror32_22_210_618;
  reg  [31:0] r8_e0_29_602;
  reg  [31:0] x_24_598;
  reg  [31:0] r1_e0_25_604;
  reg  [31:0] r4_e0_26_599;
  reg  [31:0] r6_e0_27_600;
  reg  [31:0] r3_e0_28_601;
  reg  [31:0] r2_e0_30_603;
  reg  [31:0] x_7_620;
  reg  [31:0] y_8_621;
  reg  [31:0] z_9_624;
  reg  [31:0] r3_Maj_10_627;
  reg  [31:0] r5_Maj_11_622;
  reg  [31:0] r7_Maj_12_623;
  reg  [31:0] r6_Maj_13_625;
  reg  [31:0] r4_Maj_14_626;
  reg  [31:0] arg_216_635;
  reg  [31:0] r1_ror32_6_217_639;
  reg  [5:0] r3_ror32_6_218_636;
  reg  [25:0] r6_ror32_6_219_637;
  reg  [31:0] r2_ror32_6_220_638;
  reg  [31:0] arg_176_640;
  reg  [31:0] r1_ror32_11_177_644;
  reg  [10:0] r3_ror32_11_178_641;
  reg  [20:0] r6_ror32_11_179_642;
  reg  [31:0] r2_ror32_11_180_643;
  reg  [31:0] arg_211_645;
  reg  [31:0] r1_ror32_25_212_649;
  reg  [24:0] r3_ror32_25_213_646;
  reg  [6:0] r6_ror32_25_214_647;
  reg  [31:0] r2_ror32_25_215_648;
  reg  [31:0] x_31_628;
  reg  [31:0] r1_e1_32_634;
  reg  [31:0] r4_e1_33_629;
  reg  [31:0] r6_e1_34_630;
  reg  [31:0] r3_e1_35_631;
  reg  [31:0] r8_e1_36_632;
  reg  [31:0] r2_e1_37_633;
  reg  [31:0] x_0_653;
  reg  [31:0] y_1_650;
  reg  [31:0] z_2_651;
  reg  [31:0] r3_Ch_3_656;
  reg  [31:0] r6_Ch_4_652;
  reg  [31:0] r5_Ch_5_654;
  reg  [31:0] r4_Ch_6_655;
  reg  [31:0] arg_201_664;
  reg  [31:0] r1_ror32_2_202_668;
  reg  [1:0] r3_ror32_2_203_665;
  reg  [29:0] r6_ror32_2_204_666;
  reg  [31:0] r2_ror32_2_205_667;
  reg  [31:0] arg_181_669;
  reg  [31:0] r1_ror32_13_182_673;
  reg  [12:0] r3_ror32_13_183_670;
  reg  [18:0] r6_ror32_13_184_671;
  reg  [31:0] r2_ror32_13_185_672;
  reg  [31:0] arg_206_674;
  reg  [31:0] r1_ror32_22_207_678;
  reg  [21:0] r3_ror32_22_208_675;
  reg  [9:0] r6_ror32_22_209_676;
  reg  [31:0] r2_ror32_22_210_677;
  reg  [31:0] r8_e0_29_661;
  reg  [31:0] x_24_657;
  reg  [31:0] r1_e0_25_663;
  reg  [31:0] r4_e0_26_658;
  reg  [31:0] r6_e0_27_659;
  reg  [31:0] r3_e0_28_660;
  reg  [31:0] r2_e0_30_662;
  reg  [31:0] x_7_679;
  reg  [31:0] y_8_680;
  reg  [31:0] z_9_683;
  reg  [31:0] r3_Maj_10_686;
  reg  [31:0] r5_Maj_11_681;
  reg  [31:0] r7_Maj_12_682;
  reg  [31:0] r6_Maj_13_684;
  reg  [31:0] r4_Maj_14_685;
  reg  [31:0] arg_216_694;
  reg  [31:0] r1_ror32_6_217_698;
  reg  [5:0] r3_ror32_6_218_695;
  reg  [25:0] r6_ror32_6_219_696;
  reg  [31:0] r2_ror32_6_220_697;
  reg  [31:0] arg_176_699;
  reg  [31:0] r1_ror32_11_177_703;
  reg  [10:0] r3_ror32_11_178_700;
  reg  [20:0] r6_ror32_11_179_701;
  reg  [31:0] r2_ror32_11_180_702;
  reg  [31:0] arg_211_704;
  reg  [31:0] r1_ror32_25_212_708;
  reg  [24:0] r3_ror32_25_213_705;
  reg  [6:0] r6_ror32_25_214_706;
  reg  [31:0] r2_ror32_25_215_707;
  reg  [31:0] x_31_687;
  reg  [31:0] r1_e1_32_693;
  reg  [31:0] r4_e1_33_688;
  reg  [31:0] r6_e1_34_689;
  reg  [31:0] r3_e1_35_690;
  reg  [31:0] r8_e1_36_691;
  reg  [31:0] r2_e1_37_692;
  reg  [31:0] x_0_712;
  reg  [31:0] y_1_709;
  reg  [31:0] z_2_710;
  reg  [31:0] r3_Ch_3_715;
  reg  [31:0] r6_Ch_4_711;
  reg  [31:0] r5_Ch_5_713;
  reg  [31:0] r4_Ch_6_714;
  reg  [31:0] arg_201_723;
  reg  [31:0] r1_ror32_2_202_727;
  reg  [1:0] r3_ror32_2_203_724;
  reg  [29:0] r6_ror32_2_204_725;
  reg  [31:0] r2_ror32_2_205_726;
  reg  [31:0] arg_181_728;
  reg  [31:0] r1_ror32_13_182_732;
  reg  [12:0] r3_ror32_13_183_729;
  reg  [18:0] r6_ror32_13_184_730;
  reg  [31:0] r2_ror32_13_185_731;
  reg  [31:0] arg_206_733;
  reg  [31:0] r1_ror32_22_207_737;
  reg  [21:0] r3_ror32_22_208_734;
  reg  [9:0] r6_ror32_22_209_735;
  reg  [31:0] r2_ror32_22_210_736;
  reg  [31:0] r8_e0_29_720;
  reg  [31:0] x_24_716;
  reg  [31:0] r1_e0_25_722;
  reg  [31:0] r4_e0_26_717;
  reg  [31:0] r6_e0_27_718;
  reg  [31:0] r3_e0_28_719;
  reg  [31:0] r2_e0_30_721;
  reg  [31:0] x_7_738;
  reg  [31:0] y_8_739;
  reg  [31:0] z_9_742;
  reg  [31:0] r3_Maj_10_745;
  reg  [31:0] r5_Maj_11_740;
  reg  [31:0] r7_Maj_12_741;
  reg  [31:0] r6_Maj_13_743;
  reg  [31:0] r4_Maj_14_744;
  reg  [31:0] arg_216_753;
  reg  [31:0] r1_ror32_6_217_757;
  reg  [5:0] r3_ror32_6_218_754;
  reg  [25:0] r6_ror32_6_219_755;
  reg  [31:0] r2_ror32_6_220_756;
  reg  [31:0] arg_176_758;
  reg  [31:0] r1_ror32_11_177_762;
  reg  [10:0] r3_ror32_11_178_759;
  reg  [20:0] r6_ror32_11_179_760;
  reg  [31:0] r2_ror32_11_180_761;
  reg  [31:0] arg_211_763;
  reg  [31:0] r1_ror32_25_212_767;
  reg  [24:0] r3_ror32_25_213_764;
  reg  [6:0] r6_ror32_25_214_765;
  reg  [31:0] r2_ror32_25_215_766;
  reg  [31:0] x_31_746;
  reg  [31:0] r1_e1_32_752;
  reg  [31:0] r4_e1_33_747;
  reg  [31:0] r6_e1_34_748;
  reg  [31:0] r3_e1_35_749;
  reg  [31:0] r8_e1_36_750;
  reg  [31:0] r2_e1_37_751;
  reg  [31:0] x_0_771;
  reg  [31:0] y_1_768;
  reg  [31:0] z_2_769;
  reg  [31:0] r3_Ch_3_774;
  reg  [31:0] r6_Ch_4_770;
  reg  [31:0] r5_Ch_5_772;
  reg  [31:0] r4_Ch_6_773;
  reg  [31:0] arg_201_782;
  reg  [31:0] r1_ror32_2_202_786;
  reg  [1:0] r3_ror32_2_203_783;
  reg  [29:0] r6_ror32_2_204_784;
  reg  [31:0] r2_ror32_2_205_785;
  reg  [31:0] arg_181_787;
  reg  [31:0] r1_ror32_13_182_791;
  reg  [12:0] r3_ror32_13_183_788;
  reg  [18:0] r6_ror32_13_184_789;
  reg  [31:0] r2_ror32_13_185_790;
  reg  [31:0] arg_206_792;
  reg  [31:0] r1_ror32_22_207_796;
  reg  [21:0] r3_ror32_22_208_793;
  reg  [9:0] r6_ror32_22_209_794;
  reg  [31:0] r2_ror32_22_210_795;
  reg  [31:0] r8_e0_29_779;
  reg  [31:0] x_24_775;
  reg  [31:0] r1_e0_25_781;
  reg  [31:0] r4_e0_26_776;
  reg  [31:0] r6_e0_27_777;
  reg  [31:0] r3_e0_28_778;
  reg  [31:0] r2_e0_30_780;
  reg  [31:0] x_7_797;
  reg  [31:0] y_8_798;
  reg  [31:0] z_9_801;
  reg  [31:0] r3_Maj_10_804;
  reg  [31:0] r5_Maj_11_799;
  reg  [31:0] r7_Maj_12_800;
  reg  [31:0] r6_Maj_13_802;
  reg  [31:0] r4_Maj_14_803;
  reg  [31:0] arg_216_812;
  reg  [31:0] r1_ror32_6_217_816;
  reg  [5:0] r3_ror32_6_218_813;
  reg  [25:0] r6_ror32_6_219_814;
  reg  [31:0] r2_ror32_6_220_815;
  reg  [31:0] arg_176_817;
  reg  [31:0] r1_ror32_11_177_821;
  reg  [10:0] r3_ror32_11_178_818;
  reg  [20:0] r6_ror32_11_179_819;
  reg  [31:0] r2_ror32_11_180_820;
  reg  [31:0] arg_211_822;
  reg  [31:0] r1_ror32_25_212_826;
  reg  [24:0] r3_ror32_25_213_823;
  reg  [6:0] r6_ror32_25_214_824;
  reg  [31:0] r2_ror32_25_215_825;
  reg  [31:0] x_31_805;
  reg  [31:0] r1_e1_32_811;
  reg  [31:0] r4_e1_33_806;
  reg  [31:0] r6_e1_34_807;
  reg  [31:0] r3_e1_35_808;
  reg  [31:0] r8_e1_36_809;
  reg  [31:0] r2_e1_37_810;
  reg  [31:0] x_0_830;
  reg  [31:0] y_1_827;
  reg  [31:0] z_2_828;
  reg  [31:0] r3_Ch_3_833;
  reg  [31:0] r6_Ch_4_829;
  reg  [31:0] r5_Ch_5_831;
  reg  [31:0] r4_Ch_6_832;
  reg  [31:0] arg_201_841;
  reg  [31:0] r1_ror32_2_202_845;
  reg  [1:0] r3_ror32_2_203_842;
  reg  [29:0] r6_ror32_2_204_843;
  reg  [31:0] r2_ror32_2_205_844;
  reg  [31:0] arg_181_846;
  reg  [31:0] r1_ror32_13_182_850;
  reg  [12:0] r3_ror32_13_183_847;
  reg  [18:0] r6_ror32_13_184_848;
  reg  [31:0] r2_ror32_13_185_849;
  reg  [31:0] arg_206_851;
  reg  [31:0] r1_ror32_22_207_855;
  reg  [21:0] r3_ror32_22_208_852;
  reg  [9:0] r6_ror32_22_209_853;
  reg  [31:0] r2_ror32_22_210_854;
  reg  [31:0] r8_e0_29_838;
  reg  [31:0] x_24_834;
  reg  [31:0] r1_e0_25_840;
  reg  [31:0] r4_e0_26_835;
  reg  [31:0] r6_e0_27_836;
  reg  [31:0] r3_e0_28_837;
  reg  [31:0] r2_e0_30_839;
  reg  [31:0] x_7_856;
  reg  [31:0] y_8_857;
  reg  [31:0] z_9_860;
  reg  [31:0] r3_Maj_10_863;
  reg  [31:0] r5_Maj_11_858;
  reg  [31:0] r7_Maj_12_859;
  reg  [31:0] r6_Maj_13_861;
  reg  [31:0] r4_Maj_14_862;
  reg  [31:0] arg_216_871;
  reg  [31:0] r1_ror32_6_217_875;
  reg  [5:0] r3_ror32_6_218_872;
  reg  [25:0] r6_ror32_6_219_873;
  reg  [31:0] r2_ror32_6_220_874;
  reg  [31:0] arg_176_876;
  reg  [31:0] r1_ror32_11_177_880;
  reg  [10:0] r3_ror32_11_178_877;
  reg  [20:0] r6_ror32_11_179_878;
  reg  [31:0] r2_ror32_11_180_879;
  reg  [31:0] arg_211_881;
  reg  [31:0] r1_ror32_25_212_885;
  reg  [24:0] r3_ror32_25_213_882;
  reg  [6:0] r6_ror32_25_214_883;
  reg  [31:0] r2_ror32_25_215_884;
  reg  [31:0] x_31_864;
  reg  [31:0] r1_e1_32_870;
  reg  [31:0] r4_e1_33_865;
  reg  [31:0] r6_e1_34_866;
  reg  [31:0] r3_e1_35_867;
  reg  [31:0] r8_e1_36_868;
  reg  [31:0] r2_e1_37_869;
  reg  [31:0] x_0_889;
  reg  [31:0] y_1_886;
  reg  [31:0] z_2_887;
  reg  [31:0] r3_Ch_3_892;
  reg  [31:0] r6_Ch_4_888;
  reg  [31:0] r5_Ch_5_890;
  reg  [31:0] r4_Ch_6_891;
  reg  [31:0] arg_201_900;
  reg  [31:0] r1_ror32_2_202_904;
  reg  [1:0] r3_ror32_2_203_901;
  reg  [29:0] r6_ror32_2_204_902;
  reg  [31:0] r2_ror32_2_205_903;
  reg  [31:0] arg_181_905;
  reg  [31:0] r1_ror32_13_182_909;
  reg  [12:0] r3_ror32_13_183_906;
  reg  [18:0] r6_ror32_13_184_907;
  reg  [31:0] r2_ror32_13_185_908;
  reg  [31:0] arg_206_910;
  reg  [31:0] r1_ror32_22_207_914;
  reg  [21:0] r3_ror32_22_208_911;
  reg  [9:0] r6_ror32_22_209_912;
  reg  [31:0] r2_ror32_22_210_913;
  reg  [31:0] r8_e0_29_897;
  reg  [31:0] x_24_893;
  reg  [31:0] r1_e0_25_899;
  reg  [31:0] r4_e0_26_894;
  reg  [31:0] r6_e0_27_895;
  reg  [31:0] r3_e0_28_896;
  reg  [31:0] r2_e0_30_898;
  reg  [31:0] x_7_915;
  reg  [31:0] y_8_916;
  reg  [31:0] z_9_919;
  reg  [31:0] r3_Maj_10_922;
  reg  [31:0] r5_Maj_11_917;
  reg  [31:0] r7_Maj_12_918;
  reg  [31:0] r6_Maj_13_920;
  reg  [31:0] r4_Maj_14_921;
  reg  [31:0] arg_216_930;
  reg  [31:0] r1_ror32_6_217_934;
  reg  [5:0] r3_ror32_6_218_931;
  reg  [25:0] r6_ror32_6_219_932;
  reg  [31:0] r2_ror32_6_220_933;
  reg  [31:0] arg_176_935;
  reg  [31:0] r1_ror32_11_177_939;
  reg  [10:0] r3_ror32_11_178_936;
  reg  [20:0] r6_ror32_11_179_937;
  reg  [31:0] r2_ror32_11_180_938;
  reg  [31:0] arg_211_940;
  reg  [31:0] r1_ror32_25_212_944;
  reg  [24:0] r3_ror32_25_213_941;
  reg  [6:0] r6_ror32_25_214_942;
  reg  [31:0] r2_ror32_25_215_943;
  reg  [31:0] x_31_923;
  reg  [31:0] r1_e1_32_929;
  reg  [31:0] r4_e1_33_924;
  reg  [31:0] r6_e1_34_925;
  reg  [31:0] r3_e1_35_926;
  reg  [31:0] r8_e1_36_927;
  reg  [31:0] r2_e1_37_928;
  reg  [31:0] x_0_948;
  reg  [31:0] y_1_945;
  reg  [31:0] z_2_946;
  reg  [31:0] r3_Ch_3_951;
  reg  [31:0] r6_Ch_4_947;
  reg  [31:0] r5_Ch_5_949;
  reg  [31:0] r4_Ch_6_950;
  reg  [31:0] arg_201_959;
  reg  [31:0] r1_ror32_2_202_963;
  reg  [1:0] r3_ror32_2_203_960;
  reg  [29:0] r6_ror32_2_204_961;
  reg  [31:0] r2_ror32_2_205_962;
  reg  [31:0] arg_181_964;
  reg  [31:0] r1_ror32_13_182_968;
  reg  [12:0] r3_ror32_13_183_965;
  reg  [18:0] r6_ror32_13_184_966;
  reg  [31:0] r2_ror32_13_185_967;
  reg  [31:0] arg_206_969;
  reg  [31:0] r1_ror32_22_207_973;
  reg  [21:0] r3_ror32_22_208_970;
  reg  [9:0] r6_ror32_22_209_971;
  reg  [31:0] r2_ror32_22_210_972;
  reg  [31:0] r8_e0_29_956;
  reg  [31:0] x_24_952;
  reg  [31:0] r1_e0_25_958;
  reg  [31:0] r4_e0_26_953;
  reg  [31:0] r6_e0_27_954;
  reg  [31:0] r3_e0_28_955;
  reg  [31:0] r2_e0_30_957;
  reg  [31:0] x_7_974;
  reg  [31:0] y_8_975;
  reg  [31:0] z_9_978;
  reg  [31:0] r3_Maj_10_981;
  reg  [31:0] r5_Maj_11_976;
  reg  [31:0] r7_Maj_12_977;
  reg  [31:0] r6_Maj_13_979;
  reg  [31:0] r4_Maj_14_980;
  reg  [31:0] arg_216_989;
  reg  [31:0] r1_ror32_6_217_993;
  reg  [5:0] r3_ror32_6_218_990;
  reg  [25:0] r6_ror32_6_219_991;
  reg  [31:0] r2_ror32_6_220_992;
  reg  [31:0] arg_176_994;
  reg  [31:0] r1_ror32_11_177_998;
  reg  [10:0] r3_ror32_11_178_995;
  reg  [20:0] r6_ror32_11_179_996;
  reg  [31:0] r2_ror32_11_180_997;
  reg  [31:0] arg_211_999;
  reg  [31:0] r1_ror32_25_212_1003;
  reg  [24:0] r3_ror32_25_213_1000;
  reg  [6:0] r6_ror32_25_214_1001;
  reg  [31:0] r2_ror32_25_215_1002;
  reg  [31:0] x_31_982;
  reg  [31:0] r1_e1_32_988;
  reg  [31:0] r4_e1_33_983;
  reg  [31:0] r6_e1_34_984;
  reg  [31:0] r3_e1_35_985;
  reg  [31:0] r8_e1_36_986;
  reg  [31:0] r2_e1_37_987;
  reg  [31:0] x_0_1007;
  reg  [31:0] y_1_1004;
  reg  [31:0] z_2_1005;
  reg  [31:0] r3_Ch_3_1010;
  reg  [31:0] r6_Ch_4_1006;
  reg  [31:0] r5_Ch_5_1008;
  reg  [31:0] r4_Ch_6_1009;
  reg  [31:0] arg_201_1018;
  reg  [31:0] r1_ror32_2_202_1022;
  reg  [1:0] r3_ror32_2_203_1019;
  reg  [29:0] r6_ror32_2_204_1020;
  reg  [31:0] r2_ror32_2_205_1021;
  reg  [31:0] arg_181_1023;
  reg  [31:0] r1_ror32_13_182_1027;
  reg  [12:0] r3_ror32_13_183_1024;
  reg  [18:0] r6_ror32_13_184_1025;
  reg  [31:0] r2_ror32_13_185_1026;
  reg  [31:0] arg_206_1028;
  reg  [31:0] r1_ror32_22_207_1032;
  reg  [21:0] r3_ror32_22_208_1029;
  reg  [9:0] r6_ror32_22_209_1030;
  reg  [31:0] r2_ror32_22_210_1031;
  reg  [31:0] r8_e0_29_1015;
  reg  [31:0] x_24_1011;
  reg  [31:0] r1_e0_25_1017;
  reg  [31:0] r4_e0_26_1012;
  reg  [31:0] r6_e0_27_1013;
  reg  [31:0] r3_e0_28_1014;
  reg  [31:0] r2_e0_30_1016;
  reg  [31:0] x_7_1033;
  reg  [31:0] y_8_1034;
  reg  [31:0] z_9_1037;
  reg  [31:0] r3_Maj_10_1040;
  reg  [31:0] r5_Maj_11_1035;
  reg  [31:0] r7_Maj_12_1036;
  reg  [31:0] r6_Maj_13_1038;
  reg  [31:0] r4_Maj_14_1039;
  reg  [31:0] r25_iterate_58_438;
  reg  [31:0] r78_iterate_93_478;
  reg  [31:0] r148_iterate_135_520;
  reg  [31:0] r150_iterate_136_521;
  reg  [31:0] a_39_446;
  reg  [31:0] b_40_448;
  reg  [31:0] c_41_449;
  reg  [31:0] d_42_453;
  reg  [31:0] e_43_432;
  reg  [31:0] f_44_436;
  reg  [31:0] g_45_437;
  reg  [31:0] h_46_434;
  reg  [31:0] idx_47_440;
  reg  [31:0] r9_iterate_48_561;
  reg  [31:0] r10_iterate_49_562;
  reg  [31:0] r11_iterate_50_563;
  reg  [31:0] r12_iterate_51_564;
  reg  [31:0] r13_iterate_52_565;
  reg  [31:0] r14_iterate_53_566;
  reg  [31:0] r15_iterate_54_567;
  reg  [31:0] r16_iterate_55_568;
  reg  [31:0] r23_iterate_56_433;
  reg  [31:0] r22_iterate_57_435;
  reg  [31:0] r121_iterate_118_503;
  reg  [31:0] r117_iterate_119_504;
  reg  [31:0] r21_iterate_59_439;
  reg  [31:0] r27_iterate_60_441;
  reg  [31:0] r20_iterate_61_442;
  reg  [31:0] r30_iterate_62_443;
  reg  [31:0] r19_iterate_63_444;
  reg  [31:0] r17_iterate_64_445;
  reg  [31:0] r34_iterate_65_447;
  reg  [31:0] r36_iterate_66_450;
  reg  [31:0] r33_iterate_67_451;
  reg  [31:0] r18_iterate_68_452;
  reg  [31:0] r38_iterate_69_454;
  reg  [31:0] r39_iterate_70_455;
  reg  [31:0] r44_iterate_71_456;
  reg  [31:0] r43_iterate_72_457;
  reg  [31:0] r46_iterate_73_458;
  reg  [31:0] r42_iterate_74_459;
  reg  [31:0] r48_iterate_75_460;
  reg  [31:0] r50_iterate_76_461;
  reg  [31:0] r41_iterate_77_462;
  reg  [31:0] r53_iterate_78_463;
  reg  [31:0] r55_iterate_79_464;
  reg  [31:0] r40_iterate_80_465;
  reg  [31:0] r59_iterate_81_466;
  reg  [31:0] r61_iterate_82_467;
  reg  [31:0] r58_iterate_83_468;
  reg  [31:0] r63_iterate_84_469;
  reg  [31:0] r64_iterate_85_470;
  reg  [31:0] r69_iterate_86_471;
  reg  [31:0] r68_iterate_87_472;
  reg  [31:0] r71_iterate_88_473;
  reg  [31:0] r67_iterate_89_474;
  reg  [31:0] r73_iterate_90_475;
  reg  [31:0] r75_iterate_91_476;
  reg  [31:0] r66_iterate_92_477;
  reg  [31:0] r80_iterate_94_479;
  reg  [31:0] r65_iterate_95_480;
  reg  [31:0] r84_iterate_96_481;
  reg  [31:0] r86_iterate_97_482;
  reg  [31:0] r83_iterate_98_483;
  reg  [31:0] r88_iterate_99_484;
  reg  [31:0] r89_iterate_100_485;
  reg  [31:0] r94_iterate_101_486;
  reg  [31:0] r93_iterate_102_487;
  reg  [31:0] r96_iterate_103_488;
  reg  [31:0] r92_iterate_104_489;
  reg  [31:0] r98_iterate_105_490;
  reg  [31:0] r100_iterate_106_491;
  reg  [31:0] r91_iterate_107_492;
  reg  [31:0] r103_iterate_108_493;
  reg  [31:0] r105_iterate_109_494;
  reg  [31:0] r90_iterate_110_495;
  reg  [31:0] r109_iterate_111_496;
  reg  [31:0] r111_iterate_112_497;
  reg  [31:0] r108_iterate_113_498;
  reg  [31:0] r113_iterate_114_499;
  reg  [31:0] r114_iterate_115_500;
  reg  [31:0] r213_iterate_174_559;
  reg  [31:0] r119_iterate_116_501;
  reg  [31:0] r118_iterate_117_502;
  reg  [31:0] r123_iterate_120_505;
  reg  [31:0] r125_iterate_121_506;
  reg  [31:0] r116_iterate_122_507;
  reg  [31:0] r128_iterate_123_508;
  reg  [31:0] r130_iterate_124_509;
  reg  [31:0] r115_iterate_125_510;
  reg  [31:0] r134_iterate_126_511;
  reg  [31:0] r136_iterate_127_512;
  reg  [31:0] r133_iterate_128_513;
  reg  [31:0] r138_iterate_129_514;
  reg  [31:0] r139_iterate_130_515;
  reg  [31:0] r144_iterate_131_516;
  reg  [31:0] r143_iterate_132_517;
  reg  [31:0] r146_iterate_133_518;
  reg  [31:0] r142_iterate_134_519;
  reg  [31:0] r141_iterate_137_522;
  reg  [31:0] r153_iterate_138_523;
  reg  [31:0] r155_iterate_139_524;
  reg  [31:0] r140_iterate_140_525;
  reg  [31:0] r159_iterate_141_526;
  reg  [31:0] r161_iterate_142_527;
  reg  [31:0] r158_iterate_143_528;
  reg  [31:0] r163_iterate_144_529;
  reg  [31:0] r164_iterate_145_530;
  reg  [31:0] r169_iterate_146_531;
  reg  [31:0] r168_iterate_147_532;
  reg  [31:0] r171_iterate_148_533;
  reg  [31:0] r167_iterate_149_534;
  reg  [31:0] r173_iterate_150_535;
  reg  [31:0] r175_iterate_151_536;
  reg  [31:0] r166_iterate_152_537;
  reg  [31:0] r178_iterate_153_538;
  reg  [31:0] r180_iterate_154_539;
  reg  [31:0] r165_iterate_155_540;
  reg  [31:0] r184_iterate_156_541;
  reg  [31:0] r186_iterate_157_542;
  reg  [31:0] r183_iterate_158_543;
  reg  [31:0] r188_iterate_159_544;
  reg  [31:0] r189_iterate_160_545;
  reg  [31:0] r194_iterate_161_546;
  reg  [31:0] r193_iterate_162_547;
  reg  [31:0] r196_iterate_163_548;
  reg  [31:0] r192_iterate_164_549;
  reg  [31:0] r198_iterate_165_550;
  reg  [31:0] r200_iterate_166_551;
  reg  [31:0] r191_iterate_167_552;
  reg  [31:0] r203_iterate_168_553;
  reg  [31:0] r205_iterate_169_554;
  reg  [31:0] r190_iterate_170_555;
  reg  [31:0] r209_iterate_171_556;
  reg  [31:0] r211_iterate_172_557;
  reg  [31:0] r208_iterate_173_558;
  reg  [31:0] r214_iterate_175_560;
  reg  [31:0] r__261_388;
  reg  [31:0] r0_transform_262_336;
  reg  r2_transform_263_337;
  reg  [31:0] r6_transform_264_338;
  reg  [31:0] r4_transform_265_339;
  reg  r12_transform_266_340;
  reg  [31:0] r19_transform_267_341;
  reg  [31:0] r21_transform_268_342;
  reg  [31:0] r17_transform_269_343;
  reg  [31:0] r24_transform_270_344;
  reg  [31:0] r26_transform_271_345;
  reg  [31:0] r16_transform_272_346;
  reg  [31:0] r31_transform_273_347;
  reg  [31:0] r33_transform_274_348;
  reg  [31:0] r29_transform_275_349;
  reg  [31:0] r15_transform_276_350;
  reg  [31:0] r36_transform_277_351;
  reg  [31:0] r38_transform_278_352;
  reg  [31:0] r14_transform_279_353;
  reg  [31:0] r52_transform_280_354;
  reg  [31:0] r43_transform_281_355;
  reg  [31:0] r56_transform_282_356;
  reg  [31:0] r106_transform_302_376;
  reg  [31:0] r44_transform_283_357;
  reg  [31:0] r60_transform_284_358;
  reg  [31:0] r45_transform_285_359;
  reg  [31:0] r64_transform_286_360;
  reg  [31:0] r46_transform_287_361;
  reg  [31:0] r68_transform_288_362;
  reg  [31:0] r47_transform_289_363;
  reg  [31:0] r72_transform_290_364;
  reg  [31:0] r48_transform_291_365;
  reg  [31:0] r76_transform_292_366;
  reg  [31:0] r49_transform_293_367;
  reg  [31:0] r80_transform_294_368;
  reg  [31:0] r50_transform_295_369;
  reg  r84_transform_296_370;
  reg  [31:0] r88_transform_297_371;
  reg  [31:0] r90_transform_298_372;
  reg  [31:0] r93_transform_299_373;
  reg  [31:0] r98_transform_300_374;
  reg  [31:0] r101_transform_301_375;
  reg  [31:0] r109_transform_303_377;
  reg  [31:0] r114_transform_304_378;
  reg  [31:0] r117_transform_305_379;
  reg  [31:0] r122_transform_306_380;
  reg  [31:0] r125_transform_307_381;
  reg  [31:0] r130_transform_308_382;
  reg  [31:0] r133_transform_309_383;
  reg  [31:0] r138_transform_310_384;
  reg  [31:0] r141_transform_311_385;
  reg  [31:0] r146_transform_312_386;
  reg  [31:0] r149_transform_313_387;
  reg  [31:0] addr_240_314;
  reg  [31:0] blocks_241_315;
  reg  [255:0] r2_sha256_242_334;
  reg  [31:0] r5_sha256_243_316;
  reg  r7_sha256_244_317;
  reg  [31:0] r16_sha256_245_318;
  reg  [31:0] r25_sha256_246_319;
  reg  [31:0] r29_sha256_247_320;
  reg  [63:0] r23_sha256_248_321;
  reg  [31:0] r33_sha256_249_322;
  reg  [95:0] r22_sha256_250_323;
  reg  [31:0] r37_sha256_251_324;
  reg  [127:0] r21_sha256_252_325;
  reg  [31:0] r41_sha256_253_326;
  reg  [159:0] r20_sha256_254_327;
  reg  [31:0] r45_sha256_255_328;
  reg  [191:0] r19_sha256_256_329;
  reg  [31:0] r49_sha256_257_330;
  reg  [223:0] r18_sha256_258_331;
  reg  [31:0] r53_sha256_259_332;
  reg  [255:0] r17_sha256_260_333;
  reg [31:0]  ext_task_arg_2_0;
  reg [31:0]  ext_task_arg_2_1;
  // Resources
  // add:10
  wire [31:0] add_10_s0;
  assign add_10_s0 = (st_2 == `S_2_658) ? r17_iterate_64_445 : ((st_2 == `S_2_656) ? e_43_432 : ((st_2 == `S_2_654) ? r209_iterate_171_556 : ((st_2 == `S_2_646) ? r191_iterate_167_552 : ((st_2 == `S_2_642) ? idx_47_440 : ((st_2 == `S_2_640) ? r192_iterate_164_549 : ((st_2 == `S_2_636) ? idx_47_440 : ((st_2 == `S_2_634) ? r193_iterate_162_547 : ((st_2 == `S_2_630) ? a_39_446 : ((st_2 == `S_2_625) ? r17_iterate_64_445 : ((st_2 == `S_2_623) ? f_44_436 : ((st_2 == `S_2_621) ? r184_iterate_156_541 : ((st_2 == `S_2_613) ? r166_iterate_152_537 : ((st_2 == `S_2_609) ? idx_47_440 : ((st_2 == `S_2_607) ? r167_iterate_149_534 : ((st_2 == `S_2_603) ? idx_47_440 : ((st_2 == `S_2_601) ? r168_iterate_147_532 : ((st_2 == `S_2_597) ? b_40_448 : ((st_2 == `S_2_592) ? r17_iterate_64_445 : ((st_2 == `S_2_590) ? g_45_437 : ((st_2 == `S_2_588) ? r159_iterate_141_526 : ((st_2 == `S_2_580) ? r141_iterate_137_522 : ((st_2 == `S_2_576) ? idx_47_440 : ((st_2 == `S_2_574) ? r142_iterate_134_519 : ((st_2 == `S_2_570) ? idx_47_440 : ((st_2 == `S_2_568) ? r143_iterate_132_517 : ((st_2 == `S_2_564) ? c_41_449 : ((st_2 == `S_2_559) ? r17_iterate_64_445 : ((st_2 == `S_2_557) ? h_46_434 : ((st_2 == `S_2_555) ? r134_iterate_126_511 : ((st_2 == `S_2_547) ? r116_iterate_122_507 : ((st_2 == `S_2_543) ? idx_47_440 : ((st_2 == `S_2_541) ? r117_iterate_119_504 : ((st_2 == `S_2_537) ? idx_47_440 : ((st_2 == `S_2_535) ? r118_iterate_117_502 : ((st_2 == `S_2_531) ? d_42_453 : ((st_2 == `S_2_526) ? r17_iterate_64_445 : ((st_2 == `S_2_524) ? a_39_446 : ((st_2 == `S_2_522) ? r109_iterate_111_496 : ((st_2 == `S_2_489) ? r84_iterate_96_481 : ((st_2 == `S_2_481) ? r66_iterate_92_477 : ((st_2 == `S_2_477) ? idx_47_440 : ((st_2 == `S_2_475) ? r67_iterate_89_474 : ((st_2 == `S_2_471) ? idx_47_440 : ((st_2 == `S_2_469) ? r68_iterate_87_472 : ((st_2 == `S_2_465) ? f_44_436 : ((st_2 == `S_2_460) ? r17_iterate_64_445 : ((st_2 == `S_2_458) ? c_41_449 : ((st_2 == `S_2_456) ? r59_iterate_81_466 : ((st_2 == `S_2_448) ? r41_iterate_77_462 : ((st_2 == `S_2_444) ? idx_47_440 : ((st_2 == `S_2_442) ? r42_iterate_74_459 : ((st_2 == `S_2_438) ? idx_47_440 : ((st_2 == `S_2_436) ? r43_iterate_72_457 : ((st_2 == `S_2_432) ? g_45_437 : ((st_2 == `S_2_427) ? r17_iterate_64_445 : ((st_2 == `S_2_425) ? d_42_453 : ((st_2 == `S_2_423) ? r34_iterate_65_447 : ((st_2 == `S_2_415) ? r20_iterate_61_442 : ((st_2 == `S_2_411) ? r21_iterate_59_439 : ((st_2 == `S_2_407) ? r22_iterate_57_435 : ((st_2 == `S_2_403) ? h_46_434 : ((st_2 == `S_2_286) ? r146_transform_312_386 : ((st_2 == `S_2_277) ? r138_transform_310_384 : ((st_2 == `S_2_514) ? r91_iterate_107_492 : ((st_2 == `S_2_510) ? idx_47_440 : ((st_2 == `S_2_508) ? r92_iterate_104_489 : ((st_2 == `S_2_504) ? idx_47_440 : ((st_2 == `S_2_502) ? r93_iterate_102_487 : ((st_2 == `S_2_498) ? e_43_432 : ((st_2 == `S_2_493) ? r17_iterate_64_445 : ((st_2 == `S_2_491) ? b_40_448 : ((st_2 == `S_2_241) ? r106_transform_302_376 : ((st_2 == `S_2_232) ? r98_transform_300_374 : ((st_2 == `S_2_223) ? r90_transform_298_372 : ((st_2 == `S_2_216) ? r0_transform_262_336 : ((st_2 == `S_2_165) ? r0_transform_262_336 : ((st_2 == `S_2_161) ? r15_transform_276_350 : ((st_2 == `S_2_155) ? r16_transform_272_346 : ((st_2 == `S_2_268) ? r130_transform_308_382 : ((st_2 == `S_2_259) ? r122_transform_306_380 : ((st_2 == `S_2_250) ? r114_transform_304_378 : ((st_2 == `S_2_126) ? r0_transform_262_336 : ((st_2 == `S_2_146) ? r17_transform_269_343 : ((st_2 == `S_2_21) ? r5_sha256_243_316 : (addr_240_314)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
  wire [31:0] add_10_s1;
  assign add_10_s1 = (st_2 == `S_2_658) ? r18_iterate_68_452 : ((st_2 == `S_2_656) ? r17_iterate_64_445 : ((st_2 == `S_2_654) ? r211_iterate_172_557 : ((st_2 == `S_2_646) ? r205_iterate_169_554 : ((st_2 == `S_2_642) ? 32'd7 : ((st_2 == `S_2_640) ? r200_iterate_166_551 : ((st_2 == `S_2_636) ? 32'd7 : ((st_2 == `S_2_634) ? r196_iterate_163_548 : ((st_2 == `S_2_630) ? r194_iterate_161_546 : ((st_2 == `S_2_625) ? r18_iterate_68_452 : ((st_2 == `S_2_623) ? r17_iterate_64_445 : ((st_2 == `S_2_621) ? r186_iterate_157_542 : ((st_2 == `S_2_613) ? r180_iterate_154_539 : ((st_2 == `S_2_609) ? 32'd6 : ((st_2 == `S_2_607) ? r175_iterate_151_536 : ((st_2 == `S_2_603) ? 32'd6 : ((st_2 == `S_2_601) ? r171_iterate_148_533 : ((st_2 == `S_2_597) ? r169_iterate_146_531 : ((st_2 == `S_2_592) ? r18_iterate_68_452 : ((st_2 == `S_2_590) ? r17_iterate_64_445 : ((st_2 == `S_2_588) ? r161_iterate_142_527 : ((st_2 == `S_2_580) ? r155_iterate_139_524 : ((st_2 == `S_2_576) ? 32'd5 : ((st_2 == `S_2_574) ? r150_iterate_136_521 : ((st_2 == `S_2_570) ? 32'd5 : ((st_2 == `S_2_568) ? r146_iterate_133_518 : ((st_2 == `S_2_564) ? r144_iterate_131_516 : ((st_2 == `S_2_559) ? r18_iterate_68_452 : ((st_2 == `S_2_557) ? r17_iterate_64_445 : ((st_2 == `S_2_555) ? r136_iterate_127_512 : ((st_2 == `S_2_547) ? r130_iterate_124_509 : ((st_2 == `S_2_543) ? 32'd4 : ((st_2 == `S_2_541) ? r125_iterate_121_506 : ((st_2 == `S_2_537) ? 32'd4 : ((st_2 == `S_2_535) ? r121_iterate_118_503 : ((st_2 == `S_2_531) ? r119_iterate_116_501 : ((st_2 == `S_2_526) ? r18_iterate_68_452 : ((st_2 == `S_2_524) ? r17_iterate_64_445 : ((st_2 == `S_2_522) ? r111_iterate_112_497 : ((st_2 == `S_2_489) ? r86_iterate_97_482 : ((st_2 == `S_2_481) ? r80_iterate_94_479 : ((st_2 == `S_2_477) ? 32'd2 : ((st_2 == `S_2_475) ? r75_iterate_91_476 : ((st_2 == `S_2_471) ? 32'd2 : ((st_2 == `S_2_469) ? r71_iterate_88_473 : ((st_2 == `S_2_465) ? r69_iterate_86_471 : ((st_2 == `S_2_460) ? r18_iterate_68_452 : ((st_2 == `S_2_458) ? r17_iterate_64_445 : ((st_2 == `S_2_456) ? r61_iterate_82_467 : ((st_2 == `S_2_448) ? r55_iterate_79_464 : ((st_2 == `S_2_444) ? 32'd1 : ((st_2 == `S_2_442) ? r50_iterate_76_461 : ((st_2 == `S_2_438) ? 32'd1 : ((st_2 == `S_2_436) ? r46_iterate_73_458 : ((st_2 == `S_2_432) ? r44_iterate_71_456 : ((st_2 == `S_2_427) ? r18_iterate_68_452 : ((st_2 == `S_2_425) ? r17_iterate_64_445 : ((st_2 == `S_2_423) ? r36_iterate_66_450 : ((st_2 == `S_2_415) ? r30_iterate_62_443 : ((st_2 == `S_2_411) ? r27_iterate_60_441 : ((st_2 == `S_2_407) ? r25_iterate_58_438 : ((st_2 == `S_2_403) ? r23_iterate_56_433 : ((st_2 == `S_2_286) ? r50_transform_295_369 : ((st_2 == `S_2_277) ? r49_transform_293_367 : ((st_2 == `S_2_514) ? r105_iterate_109_494 : ((st_2 == `S_2_510) ? 32'd3 : ((st_2 == `S_2_508) ? r100_iterate_106_491 : ((st_2 == `S_2_504) ? 32'd3 : ((st_2 == `S_2_502) ? r96_iterate_103_488 : ((st_2 == `S_2_498) ? r94_iterate_101_486 : ((st_2 == `S_2_493) ? r18_iterate_68_452 : ((st_2 == `S_2_491) ? r17_iterate_64_445 : ((st_2 == `S_2_241) ? r45_transform_285_359 : ((st_2 == `S_2_232) ? r44_transform_283_357 : ((st_2 == `S_2_223) ? r43_transform_281_355 : ((st_2 == `S_2_216) ? 32'd8 : ((st_2 == `S_2_165) ? 32'd1 : ((st_2 == `S_2_161) ? r38_transform_278_352 : ((st_2 == `S_2_155) ? r29_transform_275_349 : ((st_2 == `S_2_268) ? r48_transform_291_365 : ((st_2 == `S_2_259) ? r47_transform_289_363 : ((st_2 == `S_2_250) ? r46_transform_287_361 : ((st_2 == `S_2_126) ? 32'd1 : ((st_2 == `S_2_146) ? r26_transform_271_345 : ((st_2 == `S_2_21) ? 32'd1 : (32'd64)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
  wire [31:0] add_10_d0;
  assign add_10_d0 = add_10_s0 + add_10_s1;
  // gt:14
  wire [31:0] gt_14_s0;
  assign gt_14_s0 = (st_2 == `S_2_210) ? 32'd64 : ((st_2 == `S_2_131) ? 32'd64 : ((st_2 == `S_2_115) ? 32'd16 : (blocks_241_315)));
  wire [31:0] gt_14_s1;
  assign gt_14_s1 = (st_2 == `S_2_210) ? r0_transform_262_336 : ((st_2 == `S_2_131) ? r0_transform_262_336 : ((st_2 == `S_2_115) ? r0_transform_262_336 : (r5_sha256_243_316)));
  wire gt_14_d0;
  assign gt_14_d0 = gt_14_s0 > gt_14_s1;
  wire [3:0]  mem_1_2_15_p0_addr;
  wire [31:0]  mem_1_2_15_p0_rdata;
  wire [31:0]  mem_1_2_15_p0_wdata;
  wire mem_1_2_15_p0_wen;
  wire [3:0]  mem_1_2_15_p1_addr;
  wire [31:0]  mem_1_2_15_p1_rdata;
  wire [31:0]  mem_1_2_15_p1_wdata;
  wire mem_1_2_15_p1_wen;
  reg mem_1_2_15_1_2_15_ack;
  assign mem_1_2_15_p0_addr = mem_1_2_15_1_2_15_p0_addr;
  assign mem_1_2_15_p0_wdata = mem_1_2_15_1_2_15_p0_wdata;
  assign mem_1_2_15_p0_wen = (mem_1_2_15_1_2_15_p0_wen & !mem_1_2_15_1_2_15_ack);
  reg [3:0] mem_1_2_15_1_2_15_p0_addr;
  reg mem_1_2_15_1_2_15_req;
  reg [31:0] mem_1_2_15_1_2_15_p0_wdata;
  reg mem_1_2_15_1_2_15_p0_wen;
  reg [31:0] mem_1_2_15_1_2_15_rbuf;
  reg [31:0] axi_addr2_16;
  reg axi_wen2_16;
  reg axi_req2_16;
  wire axi_ack2_16;
  reg [3:0] axi_len2_16;
  reg [3:0] axi_start2_16;
  // sub:19
  wire [31:0] sub_19_s0;
  assign sub_19_s0 = (st_2 == `S_2_157) ? r0_transform_262_336 : ((st_2 == `S_2_135) ? r0_transform_262_336 : ((st_2 == `S_2_149) ? r0_transform_262_336 : (r0_transform_262_336)));
  wire [31:0] sub_19_s1;
  assign sub_19_s1 = (st_2 == `S_2_157) ? 32'd16 : ((st_2 == `S_2_135) ? 32'd2 : ((st_2 == `S_2_149) ? 32'd15 : (32'd7)));
  wire [31:0] sub_19_d0;
  assign sub_19_d0 = sub_19_s0 - sub_19_s1;
  reg [2:0] sram_addr_2;
  wire [31:0] sram_rdata_2;
  reg [31:0] sram_wdata_2;
  reg sram_wdata_en_2;
  reg [5:0] sram_addr_20;
  wire [31:0] sram_rdata_20;
  reg [31:0] sram_wdata_20;
  reg sram_wdata_en_20;
  reg [5:0] sram_addr_21;
  wire [31:0] sram_rdata_21;
  reg [31:0] sram_wdata_21;
  reg sram_wdata_en_21;
  // Insn wires
  wire  [31:0] insn_o_2_2_0;
  wire  [31:0] insn_o_2_2_1;
  wire  [31:0] insn_o_2_8_0;
  wire  insn_o_2_10_0;
  wire  [31:0] insn_o_2_25_0;
  wire  [31:0] insn_o_2_27_0;
  wire  [31:0] insn_o_2_29_0;
  wire  [31:0] insn_o_2_5_0;
  wire  [31:0] insn_o_2_14_0;
  wire  [63:0] insn_o_2_42_0;
  wire  [31:0] insn_o_2_19_0;
  wire  [95:0] insn_o_2_49_0;
  wire  [31:0] insn_o_2_22_0;
  wire  [127:0] insn_o_2_56_0;
  wire  [31:0] insn_o_2_31_0;
  wire  [159:0] insn_o_2_63_0;
  wire  [31:0] insn_o_2_35_0;
  wire  [191:0] insn_o_2_70_0;
  wire  [31:0] insn_o_2_39_0;
  wire  [223:0] insn_o_2_77_0;
  wire  [31:0] insn_o_2_45_0;
  wire  [255:0] insn_o_2_84_0;
  wire  [255:0] insn_o_2_86_0;
  wire  [31:0] insn_o_2_146_0;
  wire  insn_o_2_149_0;
  wire  [31:0] insn_o_2_155_0;
  wire  [31:0] insn_o_2_159_0;
  wire  [31:0] insn_o_2_161_0;
  wire  [31:0] insn_o_2_166_0;
  wire  [31:0] insn_o_2_170_0;
  wire  insn_o_2_173_0;
  wire  [31:0] insn_o_2_178_0;
  wire  [31:0] insn_o_2_66_0;
  wire  [31:0] insn_o_2_186_0;
  wire  [31:0] insn_o_2_188_0;
  wire  [31:0] insn_o_2_190_0;
  wire  [31:0] insn_o_2_72_0;
  wire  [31:0] insn_o_2_196_0;
  wire  [31:0] insn_o_2_200_0;
  wire  [31:0] insn_o_2_75_0;
  wire  [31:0] insn_o_2_208_0;
  wire  [31:0] insn_o_2_210_0;
  wire  [31:0] insn_o_2_211_0;
  wire  [31:0] insn_o_2_214_0;
  wire  [31:0] insn_o_2_81_0;
  wire  [31:0] insn_o_2_220_0;
  wire  [31:0] insn_o_2_226_0;
  wire  [31:0] insn_o_2_90_0;
  wire  [31:0] insn_o_2_234_0;
  wire  [31:0] insn_o_2_94_0;
  wire  [31:0] insn_o_2_241_0;
  wire  [31:0] insn_o_2_97_0;
  wire  [31:0] insn_o_2_248_0;
  wire  [31:0] insn_o_2_101_0;
  wire  [31:0] insn_o_2_255_0;
  wire  [31:0] insn_o_2_105_0;
  wire  [31:0] insn_o_2_262_0;
  wire  [31:0] insn_o_2_108_0;
  wire  [31:0] insn_o_2_269_0;
  wire  [31:0] insn_o_2_112_0;
  wire  [31:0] insn_o_2_276_0;
  wire  [31:0] insn_o_2_115_0;
  wire  [31:0] insn_o_2_283_0;
  wire  [31:0] insn_o_2_286_0;
  wire  insn_o_2_289_0;
  wire  [31:0] insn_o_2_295_0;
  wire  [31:0] insn_o_2_296_0;
  wire  [31:0] insn_o_2_297_0;
  wire  [31:0] insn_o_2_298_0;
  wire  [31:0] insn_o_2_299_0;
  wire  [31:0] insn_o_2_300_0;
  wire  [31:0] insn_o_2_301_0;
  wire  [31:0] insn_o_2_302_0;
  wire  [31:0] insn_o_2_303_0;
  wire  [31:0] insn_o_2_305_0;
  wire  [31:0] insn_o_2_306_0;
  wire  [31:0] insn_o_2_307_0;
  wire  [31:0] insn_o_2_308_0;
  wire  [31:0] insn_o_2_309_0;
  wire  [31:0] insn_o_2_310_0;
  wire  [31:0] insn_o_2_311_0;
  wire  [31:0] insn_o_2_312_0;
  wire  [31:0] insn_o_2_314_0;
  wire  [31:0] insn_o_2_316_0;
  wire  [31:0] insn_o_2_119_0;
  wire  [31:0] insn_o_2_324_0;
  wire  [31:0] insn_o_2_124_0;
  wire  [31:0] insn_o_2_336_0;
  wire  [31:0] insn_o_2_129_0;
  wire  [31:0] insn_o_2_348_0;
  wire  [31:0] insn_o_2_133_0;
  wire  [31:0] insn_o_2_360_0;
  wire  [31:0] insn_o_2_138_0;
  wire  [31:0] insn_o_2_372_0;
  wire  [31:0] insn_o_2_143_0;
  wire  [31:0] insn_o_2_384_0;
  wire  [31:0] insn_o_2_154_0;
  wire  [31:0] insn_o_2_396_0;
  wire  [31:0] insn_o_2_164_0;
  wire  [31:0] insn_o_2_408_0;
  wire  [7:0] insn_o_2_421_0;
  wire  [7:0] insn_o_2_425_0;
  wire  [15:0] insn_o_2_427_0;
  wire  [7:0] insn_o_2_431_0;
  wire  [23:0] insn_o_2_433_0;
  wire  [7:0] insn_o_2_437_0;
  wire  [31:0] insn_o_2_439_0;
  wire  [31:0] insn_o_2_441_0;
  wire  [31:0] insn_o_2_451_0;
  wire  [31:0] insn_o_2_453_0;
  wire  [31:0] insn_o_2_457_0;
  wire  [31:0] insn_o_2_459_0;
  wire  [31:0] insn_o_2_460_0;
  wire  [31:0] insn_o_2_463_0;
  wire  [31:0] insn_o_2_465_0;
  wire  [31:0] insn_o_2_467_0;
  wire  [16:0] insn_o_2_476_0;
  wire  [14:0] insn_o_2_480_0;
  wire  [31:0] insn_o_2_482_0;
  wire  [31:0] insn_o_2_484_0;
  wire  [18:0] insn_o_2_493_0;
  wire  [12:0] insn_o_2_497_0;
  wire  [31:0] insn_o_2_499_0;
  wire  [31:0] insn_o_2_501_0;
  wire  [31:0] insn_o_2_511_0;
  wire  [31:0] insn_o_2_513_0;
  wire  [31:0] insn_o_2_517_0;
  wire  [31:0] insn_o_2_519_0;
  wire  [31:0] insn_o_2_520_0;
  wire  [31:0] insn_o_2_523_0;
  wire  [31:0] insn_o_2_525_0;
  wire  [31:0] insn_o_2_527_0;
  wire  [6:0] insn_o_2_536_0;
  wire  [24:0] insn_o_2_540_0;
  wire  [31:0] insn_o_2_542_0;
  wire  [31:0] insn_o_2_544_0;
  wire  [17:0] insn_o_2_553_0;
  wire  [13:0] insn_o_2_557_0;
  wire  [31:0] insn_o_2_559_0;
  wire  [31:0] insn_o_2_561_0;
  wire  [31:0] insn_o_2_571_0;
  wire  [31:0] insn_o_2_573_0;
  wire  [31:0] insn_o_2_574_0;
  wire  [31:0] insn_o_2_579_0;
  wire  [31:0] insn_o_2_580_0;
  wire  [31:0] insn_o_2_581_0;
  wire  [31:0] insn_o_2_583_0;
  wire  [31:0] insn_o_2_584_0;
  wire  [31:0] insn_o_2_181_0;
  wire  [31:0] insn_o_2_590_0;
  wire  [31:0] insn_o_2_189_0;
  wire  [31:0] insn_o_2_596_0;
  wire  [31:0] insn_o_2_598_0;
  wire  [31:0] insn_o_2_603_0;
  wire  [31:0] insn_o_2_605_0;
  wire  [31:0] insn_o_2_609_0;
  wire  [31:0] insn_o_2_610_0;
  wire  [31:0] insn_o_2_611_0;
  wire  [31:0] insn_o_2_613_0;
  wire  [31:0] insn_o_2_614_0;
  wire  [31:0] insn_o_2_616_0;
  wire  [31:0] insn_o_2_618_0;
  wire  [31:0] insn_o_2_620_0;
  wire  [31:0] insn_o_2_622_0;
  wire  [31:0] insn_o_2_624_0;
  wire  [31:0] insn_o_2_629_0;
  wire  [31:0] insn_o_2_631_0;
  wire  [31:0] insn_o_2_632_0;
  wire  [31:0] insn_o_2_637_0;
  wire  [31:0] insn_o_2_638_0;
  wire  [31:0] insn_o_2_639_0;
  wire  [31:0] insn_o_2_641_0;
  wire  [31:0] insn_o_2_642_0;
  wire  [31:0] insn_o_2_645_0;
  wire  [31:0] insn_o_2_194_0;
  wire  [31:0] insn_o_2_651_0;
  wire  [31:0] insn_o_2_654_0;
  wire  [31:0] insn_o_2_202_0;
  wire  [31:0] insn_o_2_660_0;
  wire  [31:0] insn_o_2_662_0;
  wire  [31:0] insn_o_2_667_0;
  wire  [31:0] insn_o_2_669_0;
  wire  [31:0] insn_o_2_673_0;
  wire  [31:0] insn_o_2_674_0;
  wire  [31:0] insn_o_2_675_0;
  wire  [31:0] insn_o_2_677_0;
  wire  [31:0] insn_o_2_678_0;
  wire  [31:0] insn_o_2_680_0;
  wire  [31:0] insn_o_2_682_0;
  wire  [31:0] insn_o_2_684_0;
  wire  [31:0] insn_o_2_686_0;
  wire  [31:0] insn_o_2_688_0;
  wire  [31:0] insn_o_2_693_0;
  wire  [31:0] insn_o_2_695_0;
  wire  [31:0] insn_o_2_696_0;
  wire  [31:0] insn_o_2_701_0;
  wire  [31:0] insn_o_2_702_0;
  wire  [31:0] insn_o_2_703_0;
  wire  [31:0] insn_o_2_705_0;
  wire  [31:0] insn_o_2_706_0;
  wire  [31:0] insn_o_2_709_0;
  wire  [31:0] insn_o_2_206_0;
  wire  [31:0] insn_o_2_715_0;
  wire  [31:0] insn_o_2_718_0;
  wire  [31:0] insn_o_2_217_0;
  wire  [31:0] insn_o_2_724_0;
  wire  [31:0] insn_o_2_726_0;
  wire  [31:0] insn_o_2_731_0;
  wire  [31:0] insn_o_2_733_0;
  wire  [31:0] insn_o_2_737_0;
  wire  [31:0] insn_o_2_738_0;
  wire  [31:0] insn_o_2_739_0;
  wire  [31:0] insn_o_2_741_0;
  wire  [31:0] insn_o_2_742_0;
  wire  [31:0] insn_o_2_744_0;
  wire  [31:0] insn_o_2_746_0;
  wire  [31:0] insn_o_2_748_0;
  wire  [31:0] insn_o_2_750_0;
  wire  [31:0] insn_o_2_752_0;
  wire  [31:0] insn_o_2_757_0;
  wire  [31:0] insn_o_2_759_0;
  wire  [31:0] insn_o_2_760_0;
  wire  [31:0] insn_o_2_765_0;
  wire  [31:0] insn_o_2_766_0;
  wire  [31:0] insn_o_2_767_0;
  wire  [31:0] insn_o_2_769_0;
  wire  [31:0] insn_o_2_770_0;
  wire  [31:0] insn_o_2_773_0;
  wire  [31:0] insn_o_2_223_0;
  wire  [31:0] insn_o_2_779_0;
  wire  [31:0] insn_o_2_782_0;
  wire  [31:0] insn_o_2_230_0;
  wire  [31:0] insn_o_2_788_0;
  wire  [31:0] insn_o_2_790_0;
  wire  [31:0] insn_o_2_795_0;
  wire  [31:0] insn_o_2_797_0;
  wire  [31:0] insn_o_2_801_0;
  wire  [31:0] insn_o_2_802_0;
  wire  [31:0] insn_o_2_803_0;
  wire  [31:0] insn_o_2_805_0;
  wire  [31:0] insn_o_2_806_0;
  wire  [31:0] insn_o_2_808_0;
  wire  [31:0] insn_o_2_810_0;
  wire  [31:0] insn_o_2_812_0;
  wire  [31:0] insn_o_2_814_0;
  wire  [31:0] insn_o_2_816_0;
  wire  [31:0] insn_o_2_821_0;
  wire  [31:0] insn_o_2_823_0;
  wire  [31:0] insn_o_2_824_0;
  wire  [31:0] insn_o_2_829_0;
  wire  [31:0] insn_o_2_830_0;
  wire  [31:0] insn_o_2_831_0;
  wire  [31:0] insn_o_2_833_0;
  wire  [31:0] insn_o_2_834_0;
  wire  [31:0] insn_o_2_837_0;
  wire  [31:0] insn_o_2_236_0;
  wire  [31:0] insn_o_2_843_0;
  wire  [31:0] insn_o_2_846_0;
  wire  [31:0] insn_o_2_239_0;
  wire  [31:0] insn_o_2_852_0;
  wire  [31:0] insn_o_2_854_0;
  wire  [31:0] insn_o_2_859_0;
  wire  [31:0] insn_o_2_861_0;
  wire  [31:0] insn_o_2_865_0;
  wire  [31:0] insn_o_2_866_0;
  wire  [31:0] insn_o_2_867_0;
  wire  [31:0] insn_o_2_869_0;
  wire  [31:0] insn_o_2_870_0;
  wire  [31:0] insn_o_2_872_0;
  wire  [31:0] insn_o_2_874_0;
  wire  [31:0] insn_o_2_876_0;
  wire  [31:0] insn_o_2_878_0;
  wire  [31:0] insn_o_2_880_0;
  wire  [31:0] insn_o_2_885_0;
  wire  [31:0] insn_o_2_887_0;
  wire  [31:0] insn_o_2_888_0;
  wire  [31:0] insn_o_2_893_0;
  wire  [31:0] insn_o_2_894_0;
  wire  [31:0] insn_o_2_895_0;
  wire  [31:0] insn_o_2_897_0;
  wire  [31:0] insn_o_2_898_0;
  wire  [31:0] insn_o_2_901_0;
  wire  [31:0] insn_o_2_245_0;
  wire  [31:0] insn_o_2_907_0;
  wire  [31:0] insn_o_2_910_0;
  wire  [31:0] insn_o_2_251_0;
  wire  [31:0] insn_o_2_916_0;
  wire  [31:0] insn_o_2_918_0;
  wire  [31:0] insn_o_2_923_0;
  wire  [31:0] insn_o_2_925_0;
  wire  [31:0] insn_o_2_929_0;
  wire  [31:0] insn_o_2_930_0;
  wire  [31:0] insn_o_2_931_0;
  wire  [31:0] insn_o_2_933_0;
  wire  [31:0] insn_o_2_934_0;
  wire  [31:0] insn_o_2_936_0;
  wire  [31:0] insn_o_2_938_0;
  wire  [31:0] insn_o_2_940_0;
  wire  [31:0] insn_o_2_942_0;
  wire  [31:0] insn_o_2_944_0;
  wire  [31:0] insn_o_2_949_0;
  wire  [31:0] insn_o_2_951_0;
  wire  [31:0] insn_o_2_952_0;
  wire  [31:0] insn_o_2_957_0;
  wire  [31:0] insn_o_2_958_0;
  wire  [31:0] insn_o_2_959_0;
  wire  [31:0] insn_o_2_961_0;
  wire  [31:0] insn_o_2_962_0;
  wire  [31:0] insn_o_2_965_0;
  wire  [31:0] insn_o_2_257_0;
  wire  [31:0] insn_o_2_971_0;
  wire  [31:0] insn_o_2_974_0;
  wire  [31:0] insn_o_2_260_0;
  wire  [31:0] insn_o_2_980_0;
  wire  [31:0] insn_o_2_982_0;
  wire  [31:0] insn_o_2_987_0;
  wire  [31:0] insn_o_2_989_0;
  wire  [31:0] insn_o_2_993_0;
  wire  [31:0] insn_o_2_994_0;
  wire  [31:0] insn_o_2_995_0;
  wire  [31:0] insn_o_2_997_0;
  wire  [31:0] insn_o_2_998_0;
  wire  [31:0] insn_o_2_1000_0;
  wire  [31:0] insn_o_2_1002_0;
  wire  [31:0] insn_o_2_1004_0;
  wire  [31:0] insn_o_2_1006_0;
  wire  [31:0] insn_o_2_1008_0;
  wire  [31:0] insn_o_2_1013_0;
  wire  [31:0] insn_o_2_1015_0;
  wire  [31:0] insn_o_2_1016_0;
  wire  [31:0] insn_o_2_1021_0;
  wire  [31:0] insn_o_2_1022_0;
  wire  [31:0] insn_o_2_1023_0;
  wire  [31:0] insn_o_2_1025_0;
  wire  [31:0] insn_o_2_1026_0;
  wire  [31:0] insn_o_2_1029_0;
  wire  [31:0] insn_o_2_266_0;
  wire  [31:0] insn_o_2_1035_0;
  wire  [31:0] insn_o_2_1038_0;
  wire  [31:0] insn_o_2_272_0;
  wire  [31:0] insn_o_2_1044_0;
  wire  [31:0] insn_o_2_1046_0;
  wire  [31:0] insn_o_2_1051_0;
  wire  [31:0] insn_o_2_1053_0;
  wire  [31:0] insn_o_2_1057_0;
  wire  [31:0] insn_o_2_1058_0;
  wire  [31:0] insn_o_2_1059_0;
  wire  [31:0] insn_o_2_1061_0;
  wire  [31:0] insn_o_2_1062_0;
  wire  [31:0] insn_o_2_1064_0;
  wire  [31:0] insn_o_2_1066_0;
  wire  [31:0] insn_o_2_1068_0;
  wire  [31:0] insn_o_2_1070_0;
  wire  [31:0] insn_o_2_1072_0;
  wire  [31:0] insn_o_2_1074_0;
  wire  [31:0] insn_o_2_1076_0;
  wire  [31:0] insn_o_2_1078_0;
  wire  [31:0] insn_o_2_1080_0;
  wire  [31:0] insn_o_2_1082_0;
  wire  [31:0] insn_o_2_1084_0;
  wire  [31:0] insn_o_2_1086_0;
  wire  [31:0] insn_o_2_1088_0;
  wire  [31:0] insn_o_2_1098_0;
  wire  [31:0] insn_o_2_1100_0;
  wire  [31:0] insn_o_2_1104_0;
  wire  [31:0] insn_o_2_1106_0;
  wire  [31:0] insn_o_2_1107_0;
  wire  [31:0] insn_o_2_1112_0;
  wire  [31:0] insn_o_2_1114_0;
  wire  [31:0] insn_o_2_1115_0;
  wire  [31:0] insn_o_2_1117_0;
  wire  [5:0] insn_o_2_1126_0;
  wire  [25:0] insn_o_2_1130_0;
  wire  [31:0] insn_o_2_1132_0;
  wire  [31:0] insn_o_2_1134_0;
  wire  [10:0] insn_o_2_1143_0;
  wire  [20:0] insn_o_2_1147_0;
  wire  [31:0] insn_o_2_1149_0;
  wire  [31:0] insn_o_2_1151_0;
  wire  [24:0] insn_o_2_1160_0;
  wire  [6:0] insn_o_2_1164_0;
  wire  [31:0] insn_o_2_1166_0;
  wire  [31:0] insn_o_2_1168_0;
  wire  [31:0] insn_o_2_1175_0;
  wire  [31:0] insn_o_2_1177_0;
  wire  [31:0] insn_o_2_1179_0;
  wire  [31:0] insn_o_2_1181_0;
  wire  [31:0] insn_o_2_1191_0;
  wire  [31:0] insn_o_2_1193_0;
  wire  [31:0] insn_o_2_1197_0;
  wire  [31:0] insn_o_2_1199_0;
  wire  [31:0] insn_o_2_1200_0;
  wire  [31:0] insn_o_2_1205_0;
  wire  [31:0] insn_o_2_1207_0;
  wire  [31:0] insn_o_2_1208_0;
  wire  [31:0] insn_o_2_1210_0;
  wire  [1:0] insn_o_2_1219_0;
  wire  [29:0] insn_o_2_1223_0;
  wire  [31:0] insn_o_2_1225_0;
  wire  [31:0] insn_o_2_1227_0;
  wire  [12:0] insn_o_2_1236_0;
  wire  [18:0] insn_o_2_1240_0;
  wire  [31:0] insn_o_2_1242_0;
  wire  [31:0] insn_o_2_1244_0;
  wire  [21:0] insn_o_2_1253_0;
  wire  [9:0] insn_o_2_1257_0;
  wire  [31:0] insn_o_2_1259_0;
  wire  [31:0] insn_o_2_1261_0;
  wire  [31:0] insn_o_2_1268_0;
  wire  [31:0] insn_o_2_1270_0;
  wire  [31:0] insn_o_2_1272_0;
  wire  [31:0] insn_o_2_1274_0;
  wire  [31:0] insn_o_2_1276_0;
  wire  [31:0] insn_o_2_1286_0;
  wire  [31:0] insn_o_2_1288_0;
  wire  [31:0] insn_o_2_1292_0;
  wire  [31:0] insn_o_2_1294_0;
  wire  [31:0] insn_o_2_1295_0;
  wire  [31:0] insn_o_2_1300_0;
  wire  [31:0] insn_o_2_1302_0;
  wire  [31:0] insn_o_2_1303_0;
  wire  [31:0] insn_o_2_1305_0;
  wire  [5:0] insn_o_2_1314_0;
  wire  [25:0] insn_o_2_1318_0;
  wire  [31:0] insn_o_2_1320_0;
  wire  [31:0] insn_o_2_1322_0;
  wire  [10:0] insn_o_2_1331_0;
  wire  [20:0] insn_o_2_1335_0;
  wire  [31:0] insn_o_2_1337_0;
  wire  [31:0] insn_o_2_1339_0;
  wire  [24:0] insn_o_2_1348_0;
  wire  [6:0] insn_o_2_1352_0;
  wire  [31:0] insn_o_2_1354_0;
  wire  [31:0] insn_o_2_1356_0;
  wire  [31:0] insn_o_2_1363_0;
  wire  [31:0] insn_o_2_1365_0;
  wire  [31:0] insn_o_2_1367_0;
  wire  [31:0] insn_o_2_1369_0;
  wire  [31:0] insn_o_2_1379_0;
  wire  [31:0] insn_o_2_1381_0;
  wire  [31:0] insn_o_2_1385_0;
  wire  [31:0] insn_o_2_1387_0;
  wire  [31:0] insn_o_2_1388_0;
  wire  [31:0] insn_o_2_1393_0;
  wire  [31:0] insn_o_2_1395_0;
  wire  [31:0] insn_o_2_1396_0;
  wire  [31:0] insn_o_2_1398_0;
  wire  [1:0] insn_o_2_1407_0;
  wire  [29:0] insn_o_2_1411_0;
  wire  [31:0] insn_o_2_1413_0;
  wire  [31:0] insn_o_2_1415_0;
  wire  [12:0] insn_o_2_1424_0;
  wire  [18:0] insn_o_2_1428_0;
  wire  [31:0] insn_o_2_1430_0;
  wire  [31:0] insn_o_2_1432_0;
  wire  [21:0] insn_o_2_1441_0;
  wire  [9:0] insn_o_2_1445_0;
  wire  [31:0] insn_o_2_1447_0;
  wire  [31:0] insn_o_2_1449_0;
  wire  [31:0] insn_o_2_1456_0;
  wire  [31:0] insn_o_2_1458_0;
  wire  [31:0] insn_o_2_1460_0;
  wire  [31:0] insn_o_2_1462_0;
  wire  [31:0] insn_o_2_1464_0;
  wire  [31:0] insn_o_2_1474_0;
  wire  [31:0] insn_o_2_1476_0;
  wire  [31:0] insn_o_2_1480_0;
  wire  [31:0] insn_o_2_1482_0;
  wire  [31:0] insn_o_2_1483_0;
  wire  [31:0] insn_o_2_1488_0;
  wire  [31:0] insn_o_2_1490_0;
  wire  [31:0] insn_o_2_1491_0;
  wire  [31:0] insn_o_2_1493_0;
  wire  [5:0] insn_o_2_1502_0;
  wire  [25:0] insn_o_2_1506_0;
  wire  [31:0] insn_o_2_1508_0;
  wire  [31:0] insn_o_2_1510_0;
  wire  [10:0] insn_o_2_1519_0;
  wire  [20:0] insn_o_2_1523_0;
  wire  [31:0] insn_o_2_1525_0;
  wire  [31:0] insn_o_2_1527_0;
  wire  [24:0] insn_o_2_1536_0;
  wire  [6:0] insn_o_2_1540_0;
  wire  [31:0] insn_o_2_1542_0;
  wire  [31:0] insn_o_2_1544_0;
  wire  [31:0] insn_o_2_1551_0;
  wire  [31:0] insn_o_2_1553_0;
  wire  [31:0] insn_o_2_1555_0;
  wire  [31:0] insn_o_2_1557_0;
  wire  [31:0] insn_o_2_1567_0;
  wire  [31:0] insn_o_2_1569_0;
  wire  [31:0] insn_o_2_1573_0;
  wire  [31:0] insn_o_2_1575_0;
  wire  [31:0] insn_o_2_1576_0;
  wire  [31:0] insn_o_2_1581_0;
  wire  [31:0] insn_o_2_1583_0;
  wire  [31:0] insn_o_2_1584_0;
  wire  [31:0] insn_o_2_1586_0;
  wire  [1:0] insn_o_2_1595_0;
  wire  [29:0] insn_o_2_1599_0;
  wire  [31:0] insn_o_2_1601_0;
  wire  [31:0] insn_o_2_1603_0;
  wire  [12:0] insn_o_2_1612_0;
  wire  [18:0] insn_o_2_1616_0;
  wire  [31:0] insn_o_2_1618_0;
  wire  [31:0] insn_o_2_1620_0;
  wire  [21:0] insn_o_2_1629_0;
  wire  [9:0] insn_o_2_1633_0;
  wire  [31:0] insn_o_2_1635_0;
  wire  [31:0] insn_o_2_1637_0;
  wire  [31:0] insn_o_2_1644_0;
  wire  [31:0] insn_o_2_1646_0;
  wire  [31:0] insn_o_2_1648_0;
  wire  [31:0] insn_o_2_1650_0;
  wire  [31:0] insn_o_2_1652_0;
  wire  [31:0] insn_o_2_1662_0;
  wire  [31:0] insn_o_2_1664_0;
  wire  [31:0] insn_o_2_1668_0;
  wire  [31:0] insn_o_2_1670_0;
  wire  [31:0] insn_o_2_1671_0;
  wire  [31:0] insn_o_2_1676_0;
  wire  [31:0] insn_o_2_1678_0;
  wire  [31:0] insn_o_2_1679_0;
  wire  [31:0] insn_o_2_1681_0;
  wire  [5:0] insn_o_2_1690_0;
  wire  [25:0] insn_o_2_1694_0;
  wire  [31:0] insn_o_2_1696_0;
  wire  [31:0] insn_o_2_1698_0;
  wire  [10:0] insn_o_2_1707_0;
  wire  [20:0] insn_o_2_1711_0;
  wire  [31:0] insn_o_2_1713_0;
  wire  [31:0] insn_o_2_1715_0;
  wire  [24:0] insn_o_2_1724_0;
  wire  [6:0] insn_o_2_1728_0;
  wire  [31:0] insn_o_2_1730_0;
  wire  [31:0] insn_o_2_1732_0;
  wire  [31:0] insn_o_2_1739_0;
  wire  [31:0] insn_o_2_1741_0;
  wire  [31:0] insn_o_2_1743_0;
  wire  [31:0] insn_o_2_1745_0;
  wire  [31:0] insn_o_2_1755_0;
  wire  [31:0] insn_o_2_1757_0;
  wire  [31:0] insn_o_2_1761_0;
  wire  [31:0] insn_o_2_1763_0;
  wire  [31:0] insn_o_2_1764_0;
  wire  [31:0] insn_o_2_1769_0;
  wire  [31:0] insn_o_2_1771_0;
  wire  [31:0] insn_o_2_1772_0;
  wire  [31:0] insn_o_2_1774_0;
  wire  [1:0] insn_o_2_1783_0;
  wire  [29:0] insn_o_2_1787_0;
  wire  [31:0] insn_o_2_1789_0;
  wire  [31:0] insn_o_2_1791_0;
  wire  [12:0] insn_o_2_1800_0;
  wire  [18:0] insn_o_2_1804_0;
  wire  [31:0] insn_o_2_1806_0;
  wire  [31:0] insn_o_2_1808_0;
  wire  [21:0] insn_o_2_1817_0;
  wire  [9:0] insn_o_2_1821_0;
  wire  [31:0] insn_o_2_1823_0;
  wire  [31:0] insn_o_2_1825_0;
  wire  [31:0] insn_o_2_1832_0;
  wire  [31:0] insn_o_2_1834_0;
  wire  [31:0] insn_o_2_1836_0;
  wire  [31:0] insn_o_2_1838_0;
  wire  [31:0] insn_o_2_1840_0;
  wire  [31:0] insn_o_2_1850_0;
  wire  [31:0] insn_o_2_1852_0;
  wire  [31:0] insn_o_2_1856_0;
  wire  [31:0] insn_o_2_1858_0;
  wire  [31:0] insn_o_2_1859_0;
  wire  [31:0] insn_o_2_1864_0;
  wire  [31:0] insn_o_2_1866_0;
  wire  [31:0] insn_o_2_1867_0;
  wire  [31:0] insn_o_2_1869_0;
  wire  [5:0] insn_o_2_1878_0;
  wire  [25:0] insn_o_2_1882_0;
  wire  [31:0] insn_o_2_1884_0;
  wire  [31:0] insn_o_2_1886_0;
  wire  [10:0] insn_o_2_1895_0;
  wire  [20:0] insn_o_2_1899_0;
  wire  [31:0] insn_o_2_1901_0;
  wire  [31:0] insn_o_2_1903_0;
  wire  [24:0] insn_o_2_1912_0;
  wire  [6:0] insn_o_2_1916_0;
  wire  [31:0] insn_o_2_1918_0;
  wire  [31:0] insn_o_2_1920_0;
  wire  [31:0] insn_o_2_1927_0;
  wire  [31:0] insn_o_2_1929_0;
  wire  [31:0] insn_o_2_1931_0;
  wire  [31:0] insn_o_2_1933_0;
  wire  [31:0] insn_o_2_1943_0;
  wire  [31:0] insn_o_2_1945_0;
  wire  [31:0] insn_o_2_1949_0;
  wire  [31:0] insn_o_2_1951_0;
  wire  [31:0] insn_o_2_1952_0;
  wire  [31:0] insn_o_2_1957_0;
  wire  [31:0] insn_o_2_1959_0;
  wire  [31:0] insn_o_2_1960_0;
  wire  [31:0] insn_o_2_1962_0;
  wire  [1:0] insn_o_2_1971_0;
  wire  [29:0] insn_o_2_1975_0;
  wire  [31:0] insn_o_2_1977_0;
  wire  [31:0] insn_o_2_1979_0;
  wire  [12:0] insn_o_2_1988_0;
  wire  [18:0] insn_o_2_1992_0;
  wire  [31:0] insn_o_2_1994_0;
  wire  [31:0] insn_o_2_1996_0;
  wire  [21:0] insn_o_2_2005_0;
  wire  [9:0] insn_o_2_2009_0;
  wire  [31:0] insn_o_2_2011_0;
  wire  [31:0] insn_o_2_2013_0;
  wire  [31:0] insn_o_2_2020_0;
  wire  [31:0] insn_o_2_2022_0;
  wire  [31:0] insn_o_2_2024_0;
  wire  [31:0] insn_o_2_2026_0;
  wire  [31:0] insn_o_2_2028_0;
  wire  [31:0] insn_o_2_2038_0;
  wire  [31:0] insn_o_2_2040_0;
  wire  [31:0] insn_o_2_2044_0;
  wire  [31:0] insn_o_2_2046_0;
  wire  [31:0] insn_o_2_2047_0;
  wire  [31:0] insn_o_2_2052_0;
  wire  [31:0] insn_o_2_2054_0;
  wire  [31:0] insn_o_2_2055_0;
  wire  [31:0] insn_o_2_2057_0;
  wire  [5:0] insn_o_2_2066_0;
  wire  [25:0] insn_o_2_2070_0;
  wire  [31:0] insn_o_2_2072_0;
  wire  [31:0] insn_o_2_2074_0;
  wire  [10:0] insn_o_2_2083_0;
  wire  [20:0] insn_o_2_2087_0;
  wire  [31:0] insn_o_2_2089_0;
  wire  [31:0] insn_o_2_2091_0;
  wire  [24:0] insn_o_2_2100_0;
  wire  [6:0] insn_o_2_2104_0;
  wire  [31:0] insn_o_2_2106_0;
  wire  [31:0] insn_o_2_2108_0;
  wire  [31:0] insn_o_2_2115_0;
  wire  [31:0] insn_o_2_2117_0;
  wire  [31:0] insn_o_2_2119_0;
  wire  [31:0] insn_o_2_2121_0;
  wire  [31:0] insn_o_2_2131_0;
  wire  [31:0] insn_o_2_2133_0;
  wire  [31:0] insn_o_2_2137_0;
  wire  [31:0] insn_o_2_2139_0;
  wire  [31:0] insn_o_2_2140_0;
  wire  [31:0] insn_o_2_2145_0;
  wire  [31:0] insn_o_2_2147_0;
  wire  [31:0] insn_o_2_2148_0;
  wire  [31:0] insn_o_2_2150_0;
  wire  [1:0] insn_o_2_2159_0;
  wire  [29:0] insn_o_2_2163_0;
  wire  [31:0] insn_o_2_2165_0;
  wire  [31:0] insn_o_2_2167_0;
  wire  [12:0] insn_o_2_2176_0;
  wire  [18:0] insn_o_2_2180_0;
  wire  [31:0] insn_o_2_2182_0;
  wire  [31:0] insn_o_2_2184_0;
  wire  [21:0] insn_o_2_2193_0;
  wire  [9:0] insn_o_2_2197_0;
  wire  [31:0] insn_o_2_2199_0;
  wire  [31:0] insn_o_2_2201_0;
  wire  [31:0] insn_o_2_2208_0;
  wire  [31:0] insn_o_2_2210_0;
  wire  [31:0] insn_o_2_2212_0;
  wire  [31:0] insn_o_2_2214_0;
  wire  [31:0] insn_o_2_2216_0;
  wire  [31:0] insn_o_2_2226_0;
  wire  [31:0] insn_o_2_2228_0;
  wire  [31:0] insn_o_2_2232_0;
  wire  [31:0] insn_o_2_2234_0;
  wire  [31:0] insn_o_2_2235_0;
  wire  [31:0] insn_o_2_2240_0;
  wire  [31:0] insn_o_2_2242_0;
  wire  [31:0] insn_o_2_2243_0;
  wire  [31:0] insn_o_2_2245_0;
  wire  [5:0] insn_o_2_2254_0;
  wire  [25:0] insn_o_2_2258_0;
  wire  [31:0] insn_o_2_2260_0;
  wire  [31:0] insn_o_2_2262_0;
  wire  [10:0] insn_o_2_2271_0;
  wire  [20:0] insn_o_2_2275_0;
  wire  [31:0] insn_o_2_2277_0;
  wire  [31:0] insn_o_2_2279_0;
  wire  [24:0] insn_o_2_2288_0;
  wire  [6:0] insn_o_2_2292_0;
  wire  [31:0] insn_o_2_2294_0;
  wire  [31:0] insn_o_2_2296_0;
  wire  [31:0] insn_o_2_2303_0;
  wire  [31:0] insn_o_2_2305_0;
  wire  [31:0] insn_o_2_2307_0;
  wire  [31:0] insn_o_2_2309_0;
  wire  [31:0] insn_o_2_2319_0;
  wire  [31:0] insn_o_2_2321_0;
  wire  [31:0] insn_o_2_2325_0;
  wire  [31:0] insn_o_2_2327_0;
  wire  [31:0] insn_o_2_2328_0;
  wire  [31:0] insn_o_2_2333_0;
  wire  [31:0] insn_o_2_2335_0;
  wire  [31:0] insn_o_2_2336_0;
  wire  [31:0] insn_o_2_2338_0;
  wire  [1:0] insn_o_2_2347_0;
  wire  [29:0] insn_o_2_2351_0;
  wire  [31:0] insn_o_2_2353_0;
  wire  [31:0] insn_o_2_2355_0;
  wire  [12:0] insn_o_2_2364_0;
  wire  [18:0] insn_o_2_2368_0;
  wire  [31:0] insn_o_2_2370_0;
  wire  [31:0] insn_o_2_2372_0;
  wire  [21:0] insn_o_2_2381_0;
  wire  [9:0] insn_o_2_2385_0;
  wire  [31:0] insn_o_2_2387_0;
  wire  [31:0] insn_o_2_2389_0;
  wire  [31:0] insn_o_2_2396_0;
  wire  [31:0] insn_o_2_2398_0;
  wire  [31:0] insn_o_2_2400_0;
  wire  [31:0] insn_o_2_2402_0;
  wire  [31:0] insn_o_2_2404_0;
  wire  [31:0] insn_o_2_2414_0;
  wire  [31:0] insn_o_2_2416_0;
  wire  [31:0] insn_o_2_2420_0;
  wire  [31:0] insn_o_2_2422_0;
  wire  [31:0] insn_o_2_2423_0;
  wire  [31:0] insn_o_2_2428_0;
  wire  [31:0] insn_o_2_2430_0;
  wire  [31:0] insn_o_2_2431_0;
  wire  [31:0] insn_o_2_2433_0;
  wire  [5:0] insn_o_2_2442_0;
  wire  [25:0] insn_o_2_2446_0;
  wire  [31:0] insn_o_2_2448_0;
  wire  [31:0] insn_o_2_2450_0;
  wire  [10:0] insn_o_2_2459_0;
  wire  [20:0] insn_o_2_2463_0;
  wire  [31:0] insn_o_2_2465_0;
  wire  [31:0] insn_o_2_2467_0;
  wire  [24:0] insn_o_2_2476_0;
  wire  [6:0] insn_o_2_2480_0;
  wire  [31:0] insn_o_2_2482_0;
  wire  [31:0] insn_o_2_2484_0;
  wire  [31:0] insn_o_2_2491_0;
  wire  [31:0] insn_o_2_2493_0;
  wire  [31:0] insn_o_2_2495_0;
  wire  [31:0] insn_o_2_2497_0;
  wire  [31:0] insn_o_2_2507_0;
  wire  [31:0] insn_o_2_2509_0;
  wire  [31:0] insn_o_2_2513_0;
  wire  [31:0] insn_o_2_2515_0;
  wire  [31:0] insn_o_2_2516_0;
  wire  [31:0] insn_o_2_2521_0;
  wire  [31:0] insn_o_2_2523_0;
  wire  [31:0] insn_o_2_2524_0;
  wire  [31:0] insn_o_2_2526_0;
  wire  [1:0] insn_o_2_2535_0;
  wire  [29:0] insn_o_2_2539_0;
  wire  [31:0] insn_o_2_2541_0;
  wire  [31:0] insn_o_2_2543_0;
  wire  [12:0] insn_o_2_2552_0;
  wire  [18:0] insn_o_2_2556_0;
  wire  [31:0] insn_o_2_2558_0;
  wire  [31:0] insn_o_2_2560_0;
  wire  [21:0] insn_o_2_2569_0;
  wire  [9:0] insn_o_2_2573_0;
  wire  [31:0] insn_o_2_2575_0;
  wire  [31:0] insn_o_2_2577_0;
  wire  [31:0] insn_o_2_2584_0;
  wire  [31:0] insn_o_2_2586_0;
  wire  [31:0] insn_o_2_2588_0;
  wire  [31:0] insn_o_2_2590_0;
  wire  [31:0] insn_o_2_2592_0;
  reg [1:0] st_res_2_15;
  reg [1:0] st_res_2_16;
  reg [1:0] st_res_2_18;
  // Insn assigns
  assign insn_o_2_10_0 = gt_14_d0;
  assign insn_o_2_25_0 = add_10_d0;
  assign insn_o_2_29_0 = add_10_d0;
  assign insn_o_2_5_0 = sram_rdata_2;
  assign insn_o_2_14_0 = sram_rdata_2;
  assign insn_o_2_42_0 = {r25_sha256_246_319, r29_sha256_247_320};
  assign insn_o_2_19_0 = sram_rdata_2;
  assign insn_o_2_49_0 = {r23_sha256_248_321, r33_sha256_249_322};
  assign insn_o_2_22_0 = sram_rdata_2;
  assign insn_o_2_56_0 = {r22_sha256_250_323, r37_sha256_251_324};
  assign insn_o_2_31_0 = sram_rdata_2;
  assign insn_o_2_63_0 = {r21_sha256_252_325, r41_sha256_253_326};
  assign insn_o_2_35_0 = sram_rdata_2;
  assign insn_o_2_70_0 = {r20_sha256_254_327, r45_sha256_255_328};
  assign insn_o_2_39_0 = sram_rdata_2;
  assign insn_o_2_77_0 = {r19_sha256_256_329, r49_sha256_257_330};
  assign insn_o_2_45_0 = sram_rdata_2;
  assign insn_o_2_84_0 = {r18_sha256_258_331, r53_sha256_259_332};
  assign insn_o_2_149_0 = gt_14_d0;
  assign insn_o_2_155_0 = mem_1_2_15_1_2_15_rbuf;
  assign insn_o_2_166_0 = add_10_d0;
  assign insn_o_2_173_0 = gt_14_d0;
  assign insn_o_2_178_0 = sub_19_d0;
  assign insn_o_2_66_0 = sram_rdata_21;
  assign insn_o_2_190_0 = sub_19_d0;
  assign insn_o_2_72_0 = sram_rdata_21;
  assign insn_o_2_196_0 = add_10_d0;
  assign insn_o_2_200_0 = sub_19_d0;
  assign insn_o_2_75_0 = sram_rdata_21;
  assign insn_o_2_211_0 = add_10_d0;
  assign insn_o_2_214_0 = sub_19_d0;
  assign insn_o_2_81_0 = sram_rdata_21;
  assign insn_o_2_220_0 = add_10_d0;
  assign insn_o_2_226_0 = add_10_d0;
  assign insn_o_2_90_0 = sram_rdata_2;
  assign insn_o_2_94_0 = sram_rdata_2;
  assign insn_o_2_97_0 = sram_rdata_2;
  assign insn_o_2_101_0 = sram_rdata_2;
  assign insn_o_2_105_0 = sram_rdata_2;
  assign insn_o_2_108_0 = sram_rdata_2;
  assign insn_o_2_112_0 = sram_rdata_2;
  assign insn_o_2_115_0 = sram_rdata_2;
  assign insn_o_2_289_0 = gt_14_d0;
  assign insn_o_2_314_0 = add_10_d0;
  assign insn_o_2_119_0 = sram_rdata_2;
  assign insn_o_2_324_0 = add_10_d0;
  assign insn_o_2_124_0 = sram_rdata_2;
  assign insn_o_2_336_0 = add_10_d0;
  assign insn_o_2_129_0 = sram_rdata_2;
  assign insn_o_2_348_0 = add_10_d0;
  assign insn_o_2_133_0 = sram_rdata_2;
  assign insn_o_2_360_0 = add_10_d0;
  assign insn_o_2_138_0 = sram_rdata_2;
  assign insn_o_2_372_0 = add_10_d0;
  assign insn_o_2_143_0 = sram_rdata_2;
  assign insn_o_2_384_0 = add_10_d0;
  assign insn_o_2_154_0 = sram_rdata_2;
  assign insn_o_2_396_0 = add_10_d0;
  assign insn_o_2_164_0 = sram_rdata_2;
  assign insn_o_2_408_0 = add_10_d0;
  assign insn_o_2_421_0 = arg_15_389[7:0];
  assign insn_o_2_425_0 = arg_15_389[15:8];
  assign insn_o_2_427_0 = {r5_bswap_17_390, r8_bswap_18_391};
  assign insn_o_2_431_0 = arg_15_389[23:16];
  assign insn_o_2_433_0 = {r4_bswap_19_392, r11_bswap_20_393};
  assign insn_o_2_437_0 = arg_15_389[31:24];
  assign insn_o_2_439_0 = {r3_bswap_21_394, r14_bswap_22_395};
  assign insn_o_2_460_0 = r4_s1_235_399 ^ r6_s1_236_400;
  assign insn_o_2_463_0 = x_233_398 >> 10;
  assign insn_o_2_465_0 = r3_s1_237_401 ^ r8_s1_238_402;
  assign insn_o_2_476_0 = arg_186_405[16:0];
  assign insn_o_2_480_0 = arg_186_405[31:17];
  assign insn_o_2_482_0 = {r3_ror32_17_188_406, r6_ror32_17_189_407};
  assign insn_o_2_493_0 = arg_196_410[18:0];
  assign insn_o_2_497_0 = arg_196_410[31:19];
  assign insn_o_2_499_0 = {r3_ror32_19_198_411, r6_ror32_19_199_412};
  assign insn_o_2_520_0 = r4_s0_228_416 ^ r6_s0_229_417;
  assign insn_o_2_523_0 = x_226_415 >> 3;
  assign insn_o_2_525_0 = r3_s0_230_418 ^ r8_s0_231_419;
  assign insn_o_2_536_0 = arg_221_422[6:0];
  assign insn_o_2_540_0 = arg_221_422[31:7];
  assign insn_o_2_542_0 = {r3_ror32_7_223_423, r6_ror32_7_224_424};
  assign insn_o_2_553_0 = arg_191_427[17:0];
  assign insn_o_2_557_0 = arg_191_427[31:18];
  assign insn_o_2_559_0 = {r3_ror32_18_193_428, r6_ror32_18_194_429};
  assign insn_o_2_574_0 = add_10_d0;
  assign insn_o_2_584_0 = add_10_d0;
  assign insn_o_2_181_0 = sram_rdata_20;
  assign insn_o_2_590_0 = add_10_d0;
  assign insn_o_2_189_0 = sram_rdata_21;
  assign insn_o_2_596_0 = add_10_d0;
  assign insn_o_2_614_0 = add_10_d0;
  assign insn_o_2_618_0 = add_10_d0;
  assign insn_o_2_622_0 = add_10_d0;
  assign insn_o_2_632_0 = add_10_d0;
  assign insn_o_2_642_0 = add_10_d0;
  assign insn_o_2_645_0 = add_10_d0;
  assign insn_o_2_194_0 = sram_rdata_20;
  assign insn_o_2_651_0 = add_10_d0;
  assign insn_o_2_654_0 = add_10_d0;
  assign insn_o_2_202_0 = sram_rdata_21;
  assign insn_o_2_660_0 = add_10_d0;
  assign insn_o_2_678_0 = add_10_d0;
  assign insn_o_2_682_0 = add_10_d0;
  assign insn_o_2_686_0 = add_10_d0;
  assign insn_o_2_696_0 = add_10_d0;
  assign insn_o_2_706_0 = add_10_d0;
  assign insn_o_2_709_0 = add_10_d0;
  assign insn_o_2_206_0 = sram_rdata_20;
  assign insn_o_2_715_0 = add_10_d0;
  assign insn_o_2_718_0 = add_10_d0;
  assign insn_o_2_217_0 = sram_rdata_21;
  assign insn_o_2_724_0 = add_10_d0;
  assign insn_o_2_742_0 = add_10_d0;
  assign insn_o_2_746_0 = add_10_d0;
  assign insn_o_2_750_0 = add_10_d0;
  assign insn_o_2_760_0 = add_10_d0;
  assign insn_o_2_770_0 = add_10_d0;
  assign insn_o_2_773_0 = add_10_d0;
  assign insn_o_2_223_0 = sram_rdata_20;
  assign insn_o_2_779_0 = add_10_d0;
  assign insn_o_2_782_0 = add_10_d0;
  assign insn_o_2_230_0 = sram_rdata_21;
  assign insn_o_2_788_0 = add_10_d0;
  assign insn_o_2_806_0 = add_10_d0;
  assign insn_o_2_810_0 = add_10_d0;
  assign insn_o_2_814_0 = add_10_d0;
  assign insn_o_2_824_0 = add_10_d0;
  assign insn_o_2_834_0 = add_10_d0;
  assign insn_o_2_837_0 = add_10_d0;
  assign insn_o_2_236_0 = sram_rdata_20;
  assign insn_o_2_843_0 = add_10_d0;
  assign insn_o_2_846_0 = add_10_d0;
  assign insn_o_2_239_0 = sram_rdata_21;
  assign insn_o_2_852_0 = add_10_d0;
  assign insn_o_2_870_0 = add_10_d0;
  assign insn_o_2_874_0 = add_10_d0;
  assign insn_o_2_878_0 = add_10_d0;
  assign insn_o_2_888_0 = add_10_d0;
  assign insn_o_2_898_0 = add_10_d0;
  assign insn_o_2_901_0 = add_10_d0;
  assign insn_o_2_245_0 = sram_rdata_20;
  assign insn_o_2_907_0 = add_10_d0;
  assign insn_o_2_910_0 = add_10_d0;
  assign insn_o_2_251_0 = sram_rdata_21;
  assign insn_o_2_916_0 = add_10_d0;
  assign insn_o_2_934_0 = add_10_d0;
  assign insn_o_2_938_0 = add_10_d0;
  assign insn_o_2_942_0 = add_10_d0;
  assign insn_o_2_952_0 = add_10_d0;
  assign insn_o_2_962_0 = add_10_d0;
  assign insn_o_2_965_0 = add_10_d0;
  assign insn_o_2_257_0 = sram_rdata_20;
  assign insn_o_2_971_0 = add_10_d0;
  assign insn_o_2_974_0 = add_10_d0;
  assign insn_o_2_260_0 = sram_rdata_21;
  assign insn_o_2_980_0 = add_10_d0;
  assign insn_o_2_998_0 = add_10_d0;
  assign insn_o_2_1002_0 = add_10_d0;
  assign insn_o_2_1006_0 = add_10_d0;
  assign insn_o_2_1016_0 = add_10_d0;
  assign insn_o_2_1026_0 = add_10_d0;
  assign insn_o_2_1029_0 = add_10_d0;
  assign insn_o_2_266_0 = sram_rdata_20;
  assign insn_o_2_1035_0 = add_10_d0;
  assign insn_o_2_1038_0 = add_10_d0;
  assign insn_o_2_272_0 = sram_rdata_21;
  assign insn_o_2_1044_0 = add_10_d0;
  assign insn_o_2_1062_0 = add_10_d0;
  assign insn_o_2_1066_0 = add_10_d0;
  assign insn_o_2_1070_0 = add_10_d0;
  assign insn_o_2_1107_0 = r4_e1_33_570 ^ r6_e1_34_571;
  assign insn_o_2_1115_0 = r3_e1_35_572 ^ r8_e1_36_573;
  assign insn_o_2_1126_0 = arg_216_576[5:0];
  assign insn_o_2_1130_0 = arg_216_576[31:6];
  assign insn_o_2_1132_0 = {r3_ror32_6_218_577, r6_ror32_6_219_578};
  assign insn_o_2_1143_0 = arg_176_581[10:0];
  assign insn_o_2_1147_0 = arg_176_581[31:11];
  assign insn_o_2_1149_0 = {r3_ror32_11_178_582, r6_ror32_11_179_583};
  assign insn_o_2_1160_0 = arg_211_586[24:0];
  assign insn_o_2_1164_0 = arg_211_586[31:25];
  assign insn_o_2_1166_0 = {r3_ror32_25_213_587, r6_ror32_25_214_588};
  assign insn_o_2_1175_0 = y_1_591 ^ z_2_592;
  assign insn_o_2_1177_0 = x_0_594 & r6_Ch_4_593;
  assign insn_o_2_1179_0 = z_2_592 ^ r5_Ch_5_595;
  assign insn_o_2_1200_0 = r4_e0_26_599 ^ r6_e0_27_600;
  assign insn_o_2_1208_0 = r3_e0_28_601 ^ r8_e0_29_602;
  assign insn_o_2_1219_0 = arg_201_605[1:0];
  assign insn_o_2_1223_0 = arg_201_605[31:2];
  assign insn_o_2_1225_0 = {r3_ror32_2_203_606, r6_ror32_2_204_607};
  assign insn_o_2_1236_0 = arg_181_610[12:0];
  assign insn_o_2_1240_0 = arg_181_610[31:13];
  assign insn_o_2_1242_0 = {r3_ror32_13_183_611, r6_ror32_13_184_612};
  assign insn_o_2_1253_0 = arg_206_615[21:0];
  assign insn_o_2_1257_0 = arg_206_615[31:22];
  assign insn_o_2_1259_0 = {r3_ror32_22_208_616, r6_ror32_22_209_617};
  assign insn_o_2_1268_0 = x_7_620 & y_8_621;
  assign insn_o_2_1270_0 = x_7_620 | y_8_621;
  assign insn_o_2_1272_0 = z_9_624 & r7_Maj_12_623;
  assign insn_o_2_1274_0 = r5_Maj_11_622 | r6_Maj_13_625;
  assign insn_o_2_1295_0 = r4_e1_33_629 ^ r6_e1_34_630;
  assign insn_o_2_1303_0 = r3_e1_35_631 ^ r8_e1_36_632;
  assign insn_o_2_1314_0 = arg_216_635[5:0];
  assign insn_o_2_1318_0 = arg_216_635[31:6];
  assign insn_o_2_1320_0 = {r3_ror32_6_218_636, r6_ror32_6_219_637};
  assign insn_o_2_1331_0 = arg_176_640[10:0];
  assign insn_o_2_1335_0 = arg_176_640[31:11];
  assign insn_o_2_1337_0 = {r3_ror32_11_178_641, r6_ror32_11_179_642};
  assign insn_o_2_1348_0 = arg_211_645[24:0];
  assign insn_o_2_1352_0 = arg_211_645[31:25];
  assign insn_o_2_1354_0 = {r3_ror32_25_213_646, r6_ror32_25_214_647};
  assign insn_o_2_1363_0 = y_1_650 ^ z_2_651;
  assign insn_o_2_1365_0 = x_0_653 & r6_Ch_4_652;
  assign insn_o_2_1367_0 = z_2_651 ^ r5_Ch_5_654;
  assign insn_o_2_1388_0 = r4_e0_26_658 ^ r6_e0_27_659;
  assign insn_o_2_1396_0 = r3_e0_28_660 ^ r8_e0_29_661;
  assign insn_o_2_1407_0 = arg_201_664[1:0];
  assign insn_o_2_1411_0 = arg_201_664[31:2];
  assign insn_o_2_1413_0 = {r3_ror32_2_203_665, r6_ror32_2_204_666};
  assign insn_o_2_1424_0 = arg_181_669[12:0];
  assign insn_o_2_1428_0 = arg_181_669[31:13];
  assign insn_o_2_1430_0 = {r3_ror32_13_183_670, r6_ror32_13_184_671};
  assign insn_o_2_1441_0 = arg_206_674[21:0];
  assign insn_o_2_1445_0 = arg_206_674[31:22];
  assign insn_o_2_1447_0 = {r3_ror32_22_208_675, r6_ror32_22_209_676};
  assign insn_o_2_1456_0 = x_7_679 & y_8_680;
  assign insn_o_2_1458_0 = x_7_679 | y_8_680;
  assign insn_o_2_1460_0 = z_9_683 & r7_Maj_12_682;
  assign insn_o_2_1462_0 = r5_Maj_11_681 | r6_Maj_13_684;
  assign insn_o_2_1483_0 = r4_e1_33_688 ^ r6_e1_34_689;
  assign insn_o_2_1491_0 = r3_e1_35_690 ^ r8_e1_36_691;
  assign insn_o_2_1502_0 = arg_216_694[5:0];
  assign insn_o_2_1506_0 = arg_216_694[31:6];
  assign insn_o_2_1508_0 = {r3_ror32_6_218_695, r6_ror32_6_219_696};
  assign insn_o_2_1519_0 = arg_176_699[10:0];
  assign insn_o_2_1523_0 = arg_176_699[31:11];
  assign insn_o_2_1525_0 = {r3_ror32_11_178_700, r6_ror32_11_179_701};
  assign insn_o_2_1536_0 = arg_211_704[24:0];
  assign insn_o_2_1540_0 = arg_211_704[31:25];
  assign insn_o_2_1542_0 = {r3_ror32_25_213_705, r6_ror32_25_214_706};
  assign insn_o_2_1551_0 = y_1_709 ^ z_2_710;
  assign insn_o_2_1553_0 = x_0_712 & r6_Ch_4_711;
  assign insn_o_2_1555_0 = z_2_710 ^ r5_Ch_5_713;
  assign insn_o_2_1576_0 = r4_e0_26_717 ^ r6_e0_27_718;
  assign insn_o_2_1584_0 = r3_e0_28_719 ^ r8_e0_29_720;
  assign insn_o_2_1595_0 = arg_201_723[1:0];
  assign insn_o_2_1599_0 = arg_201_723[31:2];
  assign insn_o_2_1601_0 = {r3_ror32_2_203_724, r6_ror32_2_204_725};
  assign insn_o_2_1612_0 = arg_181_728[12:0];
  assign insn_o_2_1616_0 = arg_181_728[31:13];
  assign insn_o_2_1618_0 = {r3_ror32_13_183_729, r6_ror32_13_184_730};
  assign insn_o_2_1629_0 = arg_206_733[21:0];
  assign insn_o_2_1633_0 = arg_206_733[31:22];
  assign insn_o_2_1635_0 = {r3_ror32_22_208_734, r6_ror32_22_209_735};
  assign insn_o_2_1644_0 = x_7_738 & y_8_739;
  assign insn_o_2_1646_0 = x_7_738 | y_8_739;
  assign insn_o_2_1648_0 = z_9_742 & r7_Maj_12_741;
  assign insn_o_2_1650_0 = r5_Maj_11_740 | r6_Maj_13_743;
  assign insn_o_2_1671_0 = r4_e1_33_747 ^ r6_e1_34_748;
  assign insn_o_2_1679_0 = r3_e1_35_749 ^ r8_e1_36_750;
  assign insn_o_2_1690_0 = arg_216_753[5:0];
  assign insn_o_2_1694_0 = arg_216_753[31:6];
  assign insn_o_2_1696_0 = {r3_ror32_6_218_754, r6_ror32_6_219_755};
  assign insn_o_2_1707_0 = arg_176_758[10:0];
  assign insn_o_2_1711_0 = arg_176_758[31:11];
  assign insn_o_2_1713_0 = {r3_ror32_11_178_759, r6_ror32_11_179_760};
  assign insn_o_2_1724_0 = arg_211_763[24:0];
  assign insn_o_2_1728_0 = arg_211_763[31:25];
  assign insn_o_2_1730_0 = {r3_ror32_25_213_764, r6_ror32_25_214_765};
  assign insn_o_2_1739_0 = y_1_768 ^ z_2_769;
  assign insn_o_2_1741_0 = x_0_771 & r6_Ch_4_770;
  assign insn_o_2_1743_0 = z_2_769 ^ r5_Ch_5_772;
  assign insn_o_2_1764_0 = r4_e0_26_776 ^ r6_e0_27_777;
  assign insn_o_2_1772_0 = r3_e0_28_778 ^ r8_e0_29_779;
  assign insn_o_2_1783_0 = arg_201_782[1:0];
  assign insn_o_2_1787_0 = arg_201_782[31:2];
  assign insn_o_2_1789_0 = {r3_ror32_2_203_783, r6_ror32_2_204_784};
  assign insn_o_2_1800_0 = arg_181_787[12:0];
  assign insn_o_2_1804_0 = arg_181_787[31:13];
  assign insn_o_2_1806_0 = {r3_ror32_13_183_788, r6_ror32_13_184_789};
  assign insn_o_2_1817_0 = arg_206_792[21:0];
  assign insn_o_2_1821_0 = arg_206_792[31:22];
  assign insn_o_2_1823_0 = {r3_ror32_22_208_793, r6_ror32_22_209_794};
  assign insn_o_2_1832_0 = x_7_797 & y_8_798;
  assign insn_o_2_1834_0 = x_7_797 | y_8_798;
  assign insn_o_2_1836_0 = z_9_801 & r7_Maj_12_800;
  assign insn_o_2_1838_0 = r5_Maj_11_799 | r6_Maj_13_802;
  assign insn_o_2_1859_0 = r4_e1_33_806 ^ r6_e1_34_807;
  assign insn_o_2_1867_0 = r3_e1_35_808 ^ r8_e1_36_809;
  assign insn_o_2_1878_0 = arg_216_812[5:0];
  assign insn_o_2_1882_0 = arg_216_812[31:6];
  assign insn_o_2_1884_0 = {r3_ror32_6_218_813, r6_ror32_6_219_814};
  assign insn_o_2_1895_0 = arg_176_817[10:0];
  assign insn_o_2_1899_0 = arg_176_817[31:11];
  assign insn_o_2_1901_0 = {r3_ror32_11_178_818, r6_ror32_11_179_819};
  assign insn_o_2_1912_0 = arg_211_822[24:0];
  assign insn_o_2_1916_0 = arg_211_822[31:25];
  assign insn_o_2_1918_0 = {r3_ror32_25_213_823, r6_ror32_25_214_824};
  assign insn_o_2_1927_0 = y_1_827 ^ z_2_828;
  assign insn_o_2_1929_0 = x_0_830 & r6_Ch_4_829;
  assign insn_o_2_1931_0 = z_2_828 ^ r5_Ch_5_831;
  assign insn_o_2_1952_0 = r4_e0_26_835 ^ r6_e0_27_836;
  assign insn_o_2_1960_0 = r3_e0_28_837 ^ r8_e0_29_838;
  assign insn_o_2_1971_0 = arg_201_841[1:0];
  assign insn_o_2_1975_0 = arg_201_841[31:2];
  assign insn_o_2_1977_0 = {r3_ror32_2_203_842, r6_ror32_2_204_843};
  assign insn_o_2_1988_0 = arg_181_846[12:0];
  assign insn_o_2_1992_0 = arg_181_846[31:13];
  assign insn_o_2_1994_0 = {r3_ror32_13_183_847, r6_ror32_13_184_848};
  assign insn_o_2_2005_0 = arg_206_851[21:0];
  assign insn_o_2_2009_0 = arg_206_851[31:22];
  assign insn_o_2_2011_0 = {r3_ror32_22_208_852, r6_ror32_22_209_853};
  assign insn_o_2_2020_0 = x_7_856 & y_8_857;
  assign insn_o_2_2022_0 = x_7_856 | y_8_857;
  assign insn_o_2_2024_0 = z_9_860 & r7_Maj_12_859;
  assign insn_o_2_2026_0 = r5_Maj_11_858 | r6_Maj_13_861;
  assign insn_o_2_2047_0 = r4_e1_33_865 ^ r6_e1_34_866;
  assign insn_o_2_2055_0 = r3_e1_35_867 ^ r8_e1_36_868;
  assign insn_o_2_2066_0 = arg_216_871[5:0];
  assign insn_o_2_2070_0 = arg_216_871[31:6];
  assign insn_o_2_2072_0 = {r3_ror32_6_218_872, r6_ror32_6_219_873};
  assign insn_o_2_2083_0 = arg_176_876[10:0];
  assign insn_o_2_2087_0 = arg_176_876[31:11];
  assign insn_o_2_2089_0 = {r3_ror32_11_178_877, r6_ror32_11_179_878};
  assign insn_o_2_2100_0 = arg_211_881[24:0];
  assign insn_o_2_2104_0 = arg_211_881[31:25];
  assign insn_o_2_2106_0 = {r3_ror32_25_213_882, r6_ror32_25_214_883};
  assign insn_o_2_2115_0 = y_1_886 ^ z_2_887;
  assign insn_o_2_2117_0 = x_0_889 & r6_Ch_4_888;
  assign insn_o_2_2119_0 = z_2_887 ^ r5_Ch_5_890;
  assign insn_o_2_2140_0 = r4_e0_26_894 ^ r6_e0_27_895;
  assign insn_o_2_2148_0 = r3_e0_28_896 ^ r8_e0_29_897;
  assign insn_o_2_2159_0 = arg_201_900[1:0];
  assign insn_o_2_2163_0 = arg_201_900[31:2];
  assign insn_o_2_2165_0 = {r3_ror32_2_203_901, r6_ror32_2_204_902};
  assign insn_o_2_2176_0 = arg_181_905[12:0];
  assign insn_o_2_2180_0 = arg_181_905[31:13];
  assign insn_o_2_2182_0 = {r3_ror32_13_183_906, r6_ror32_13_184_907};
  assign insn_o_2_2193_0 = arg_206_910[21:0];
  assign insn_o_2_2197_0 = arg_206_910[31:22];
  assign insn_o_2_2199_0 = {r3_ror32_22_208_911, r6_ror32_22_209_912};
  assign insn_o_2_2208_0 = x_7_915 & y_8_916;
  assign insn_o_2_2210_0 = x_7_915 | y_8_916;
  assign insn_o_2_2212_0 = z_9_919 & r7_Maj_12_918;
  assign insn_o_2_2214_0 = r5_Maj_11_917 | r6_Maj_13_920;
  assign insn_o_2_2235_0 = r4_e1_33_924 ^ r6_e1_34_925;
  assign insn_o_2_2243_0 = r3_e1_35_926 ^ r8_e1_36_927;
  assign insn_o_2_2254_0 = arg_216_930[5:0];
  assign insn_o_2_2258_0 = arg_216_930[31:6];
  assign insn_o_2_2260_0 = {r3_ror32_6_218_931, r6_ror32_6_219_932};
  assign insn_o_2_2271_0 = arg_176_935[10:0];
  assign insn_o_2_2275_0 = arg_176_935[31:11];
  assign insn_o_2_2277_0 = {r3_ror32_11_178_936, r6_ror32_11_179_937};
  assign insn_o_2_2288_0 = arg_211_940[24:0];
  assign insn_o_2_2292_0 = arg_211_940[31:25];
  assign insn_o_2_2294_0 = {r3_ror32_25_213_941, r6_ror32_25_214_942};
  assign insn_o_2_2303_0 = y_1_945 ^ z_2_946;
  assign insn_o_2_2305_0 = x_0_948 & r6_Ch_4_947;
  assign insn_o_2_2307_0 = z_2_946 ^ r5_Ch_5_949;
  assign insn_o_2_2328_0 = r4_e0_26_953 ^ r6_e0_27_954;
  assign insn_o_2_2336_0 = r3_e0_28_955 ^ r8_e0_29_956;
  assign insn_o_2_2347_0 = arg_201_959[1:0];
  assign insn_o_2_2351_0 = arg_201_959[31:2];
  assign insn_o_2_2353_0 = {r3_ror32_2_203_960, r6_ror32_2_204_961};
  assign insn_o_2_2364_0 = arg_181_964[12:0];
  assign insn_o_2_2368_0 = arg_181_964[31:13];
  assign insn_o_2_2370_0 = {r3_ror32_13_183_965, r6_ror32_13_184_966};
  assign insn_o_2_2381_0 = arg_206_969[21:0];
  assign insn_o_2_2385_0 = arg_206_969[31:22];
  assign insn_o_2_2387_0 = {r3_ror32_22_208_970, r6_ror32_22_209_971};
  assign insn_o_2_2396_0 = x_7_974 & y_8_975;
  assign insn_o_2_2398_0 = x_7_974 | y_8_975;
  assign insn_o_2_2400_0 = z_9_978 & r7_Maj_12_977;
  assign insn_o_2_2402_0 = r5_Maj_11_976 | r6_Maj_13_979;
  assign insn_o_2_2423_0 = r4_e1_33_983 ^ r6_e1_34_984;
  assign insn_o_2_2431_0 = r3_e1_35_985 ^ r8_e1_36_986;
  assign insn_o_2_2442_0 = arg_216_989[5:0];
  assign insn_o_2_2446_0 = arg_216_989[31:6];
  assign insn_o_2_2448_0 = {r3_ror32_6_218_990, r6_ror32_6_219_991};
  assign insn_o_2_2459_0 = arg_176_994[10:0];
  assign insn_o_2_2463_0 = arg_176_994[31:11];
  assign insn_o_2_2465_0 = {r3_ror32_11_178_995, r6_ror32_11_179_996};
  assign insn_o_2_2476_0 = arg_211_999[24:0];
  assign insn_o_2_2480_0 = arg_211_999[31:25];
  assign insn_o_2_2482_0 = {r3_ror32_25_213_1000, r6_ror32_25_214_1001};
  assign insn_o_2_2491_0 = y_1_1004 ^ z_2_1005;
  assign insn_o_2_2493_0 = x_0_1007 & r6_Ch_4_1006;
  assign insn_o_2_2495_0 = z_2_1005 ^ r5_Ch_5_1008;
  assign insn_o_2_2516_0 = r4_e0_26_1012 ^ r6_e0_27_1013;
  assign insn_o_2_2524_0 = r3_e0_28_1014 ^ r8_e0_29_1015;
  assign insn_o_2_2535_0 = arg_201_1018[1:0];
  assign insn_o_2_2539_0 = arg_201_1018[31:2];
  assign insn_o_2_2541_0 = {r3_ror32_2_203_1019, r6_ror32_2_204_1020};
  assign insn_o_2_2552_0 = arg_181_1023[12:0];
  assign insn_o_2_2556_0 = arg_181_1023[31:13];
  assign insn_o_2_2558_0 = {r3_ror32_13_183_1024, r6_ror32_13_184_1025};
  assign insn_o_2_2569_0 = arg_206_1028[21:0];
  assign insn_o_2_2573_0 = arg_206_1028[31:22];
  assign insn_o_2_2575_0 = {r3_ror32_22_208_1029, r6_ror32_22_209_1030};
  assign insn_o_2_2584_0 = x_7_1033 & y_8_1034;
  assign insn_o_2_2586_0 = x_7_1033 | y_8_1034;
  assign insn_o_2_2588_0 = z_9_1037 & r7_Maj_12_1036;
  assign insn_o_2_2590_0 = r5_Maj_11_1035 | r6_Maj_13_1038;
  assign insn_o_2_2_0 = ext_task_arg_2_0;
  assign insn_o_2_2_1 = ext_task_arg_2_1;

  // Table 1
  always @(posedge clk) begin
    if (rst) begin
      st_1 <= `S_1_1;
    end else begin
      case (st_1)
        `S_1_1: begin
          st_1 <= `S_1_2;
        end
        `S_1_2: begin
        end
      endcase
    end
  end
  // Table 2
  always @(posedge clk) begin
    if (rst) begin
      st_2 <= `S_2_task_idle;
      mem_1_2_15_1_2_15_ack <= 0;
      mem_1_2_15_1_2_15_req <= 0;
      mem_1_2_15_1_2_15_p0_wen <= 0;
      axi_addr2_16 <= 0;
      axi_wen2_16 <= 0;
      axi_req2_16 <= 0;
      sha256_req_ready <= 0;
      sha256_res_valid <= 0;
      sha256_req_busy <= 0;
      st_res_2_15 <= 0;
      st_res_2_16 <= 0;
      st_res_2_18 <= 0;
    end else begin
      mem_1_2_15_1_2_15_ack <= !(0) && mem_1_2_15_1_2_15_req;
      mem_1_2_15_1_2_15_req <= ((st_2 == `S_2_120 && st_res_2_15 == 0)) && !mem_1_2_15_1_2_15_ack;
      mem_1_2_15_1_2_15_p0_wen <= 0 && !mem_1_2_15_1_2_15_ack;
      axi_req2_16 <= ((st_2 == `S_2_13 && st_res_2_16 == 0)) && !axi_ack2_16;
      axi_wen2_16 <= 0;
      sha256_req_ready <= sha256_req_valid & (st_2 == `S_2_task_idle);
      sha256_req_busy <= !(st_2 == `S_2_task_idle);
      sram_wdata_en_2 <= (st_2 == 72) | (st_2 == 77) | (st_2 == 82) | (st_2 == 87) | (st_2 == 92) | (st_2 == 97) | (st_2 == 102) | (st_2 == 107) | (st_2 == 254) | (st_2 == 263) | (st_2 == 227) | (st_2 == 236) | (st_2 == 245) | (st_2 == 272) | (st_2 == 281) | (st_2 == 290);
      sram_wdata_en_20 <= 0;
      sram_wdata_en_21 <= (st_2 == 125) | (st_2 == 164);
      case (st_2)
        `S_2_task_idle: begin
          if (sha256_req_valid) begin
            st_2 <= `S_2_1;
            ext_task_arg_2_0 <= sha256_req_0;
            ext_task_arg_2_1 <= sha256_req_1;
          end
        end
        `S_2_1: begin
          addr_240_314 <= insn_o_2_2_0;
          blocks_241_315 <= insn_o_2_2_1;
          st_2 <= `S_2_72;
        end
        `S_2_6: begin
          r5_sha256_243_316 <= 32'd0;
          st_2 <= `S_2_7;
        end
        `S_2_7: begin
          r7_sha256_244_317 <= insn_o_2_10_0;
          st_2 <= `S_2_8;
        end
        `S_2_8: begin
          if (r7_sha256_244_317) begin
            st_2 <= `S_2_9;
          end else begin
            st_2 <= `S_2_23;
          end
        end
        `S_2_9: begin
          st_2 <= `S_2_13;
        end
        `S_2_13: begin
          // AXI access request
          if (st_res_2_16 == 0) begin
            axi_addr2_16 <= addr_240_314;
            axi_len2_16 <= 32'd15;
            axi_start2_16 <= 32'd0;
            if (axi_ack2_16) begin
              st_res_2_16 <= 3;
            end
          end
          if ((st_res_2_16 == 3)) begin
            // 1 cycle insns
          end
          if ((st_res_2_16 == 3)) begin
            // clears sub states
            st_res_2_16 <= 0;
          end
          if ((st_res_2_16 == 3)) begin
          st_2 <= `S_2_113;
          end
        end
        `S_2_19: begin
          r16_sha256_245_318 <= insn_o_2_25_0;
          st_2 <= `S_2_20;
        end
        `S_2_20: begin
          addr_240_314 <= r16_sha256_245_318;
          st_2 <= `S_2_21;
        end
        `S_2_21: begin
          r5_sha256_243_316 <= insn_o_2_29_0;
          st_2 <= `S_2_7;
        end
        `S_2_23: begin
          st_2 <= `S_2_26;
        end
        `S_2_26: begin
          sram_addr_2 <= 32'd0;
          st_2 <= `S_2_2;
        end
        `S_2_2: begin
          r25_sha256_246_319 <= insn_o_2_5_0;
          st_2 <= `S_2_30;
        end
        `S_2_30: begin
          sram_addr_2 <= 32'd1;
          st_2 <= `S_2_3;
        end
        `S_2_3: begin
          r29_sha256_247_320 <= insn_o_2_14_0;
          st_2 <= `S_2_31;
        end
        `S_2_31: begin
          r23_sha256_248_321 <= insn_o_2_42_0;
          st_2 <= `S_2_35;
        end
        `S_2_35: begin
          sram_addr_2 <= 32'd2;
          st_2 <= `S_2_4;
        end
        `S_2_4: begin
          r33_sha256_249_322 <= insn_o_2_19_0;
          st_2 <= `S_2_36;
        end
        `S_2_36: begin
          r22_sha256_250_323 <= insn_o_2_49_0;
          st_2 <= `S_2_40;
        end
        `S_2_40: begin
          sram_addr_2 <= 32'd3;
          st_2 <= `S_2_5;
        end
        `S_2_5: begin
          r37_sha256_251_324 <= insn_o_2_22_0;
          st_2 <= `S_2_41;
        end
        `S_2_41: begin
          r21_sha256_252_325 <= insn_o_2_56_0;
          st_2 <= `S_2_45;
        end
        `S_2_45: begin
          sram_addr_2 <= 32'd4;
          st_2 <= `S_2_10;
        end
        `S_2_10: begin
          r41_sha256_253_326 <= insn_o_2_31_0;
          st_2 <= `S_2_46;
        end
        `S_2_46: begin
          r20_sha256_254_327 <= insn_o_2_63_0;
          st_2 <= `S_2_50;
        end
        `S_2_50: begin
          sram_addr_2 <= 32'd5;
          st_2 <= `S_2_11;
        end
        `S_2_11: begin
          r45_sha256_255_328 <= insn_o_2_35_0;
          st_2 <= `S_2_51;
        end
        `S_2_51: begin
          r19_sha256_256_329 <= insn_o_2_70_0;
          st_2 <= `S_2_55;
        end
        `S_2_55: begin
          sram_addr_2 <= 32'd6;
          st_2 <= `S_2_12;
        end
        `S_2_12: begin
          r49_sha256_257_330 <= insn_o_2_39_0;
          st_2 <= `S_2_56;
        end
        `S_2_56: begin
          r18_sha256_258_331 <= insn_o_2_77_0;
          st_2 <= `S_2_60;
        end
        `S_2_60: begin
          sram_addr_2 <= 32'd7;
          st_2 <= `S_2_14;
        end
        `S_2_14: begin
          r53_sha256_259_332 <= insn_o_2_45_0;
          st_2 <= `S_2_61;
        end
        `S_2_61: begin
          r17_sha256_260_333 <= insn_o_2_84_0;
          st_2 <= `S_2_62;
        end
        `S_2_62: begin
          r2_sha256_242_334 <= r17_sha256_260_333;
          st_2 <= `S_2_66;
        end
        `S_2_66: begin
          if (st_res_2_18 == 0) begin
            sha256_res_valid <= 1;
            st_res_2_18 <= 1;
            sha256_res_0 <= r2_sha256_242_334;
          end
          if (st_res_2_18 == 1) begin
            if (sha256_res_ready) begin
              sha256_res_valid <= 0;
              st_res_2_18 <= 3;
            end
          end
          if ((st_res_2_18 == 3)) begin
            // 1 cycle insns
          end
          if ((st_res_2_18 == 3)) begin
            // clears sub states
            st_res_2_18 <= 0;
          end
          if ((st_res_2_18 == 3)) begin
          st_2 <= `S_2_task_idle;
          end
        end
        `S_2_72: begin
          sram_addr_2 <= 32'd0;
          sram_wdata_2 <= 32'd1779033703;
          st_2 <= `S_2_77;
        end
        `S_2_77: begin
          sram_addr_2 <= 32'd1;
          sram_wdata_2 <= 32'd2147483647;
          st_2 <= `S_2_82;
        end
        `S_2_82: begin
          sram_addr_2 <= 32'd2;
          sram_wdata_2 <= 32'd1013904242;
          st_2 <= `S_2_87;
        end
        `S_2_87: begin
          sram_addr_2 <= 32'd3;
          sram_wdata_2 <= 32'd2147483647;
          st_2 <= `S_2_92;
        end
        `S_2_92: begin
          sram_addr_2 <= 32'd4;
          sram_wdata_2 <= 32'd1359893119;
          st_2 <= `S_2_97;
        end
        `S_2_97: begin
          sram_addr_2 <= 32'd5;
          sram_wdata_2 <= 32'd2147483647;
          st_2 <= `S_2_102;
        end
        `S_2_102: begin
          sram_addr_2 <= 32'd6;
          sram_wdata_2 <= 32'd528734635;
          st_2 <= `S_2_107;
        end
        `S_2_107: begin
          sram_addr_2 <= 32'd7;
          sram_wdata_2 <= 32'd1541459225;
          st_2 <= `S_2_6;
        end
        `S_2_113: begin
          r0_transform_262_336 <= 32'd0;
          st_2 <= `S_2_114;
        end
        `S_2_114: begin
          st_2 <= `S_2_115;
        end
        `S_2_115: begin
          r2_transform_263_337 <= insn_o_2_149_0;
          st_2 <= `S_2_116;
        end
        `S_2_116: begin
          if (r2_transform_263_337) begin
            st_2 <= `S_2_117;
          end else begin
            st_2 <= `S_2_128;
          end
        end
        `S_2_117: begin
          st_2 <= `S_2_120;
        end
        `S_2_120: begin
          if (st_res_2_15 == 0) begin
            mem_1_2_15_1_2_15_p0_addr <= r0_transform_262_336;
            if (mem_1_2_15_1_2_15_ack) begin
              st_res_2_15 <= 3;
              mem_1_2_15_1_2_15_rbuf <= mem_1_2_15_p0_rdata;
            end
          end
          if ((st_res_2_15 == 3)) begin
            // 1 cycle insns
          r6_transform_264_338 <= insn_o_2_155_0;
          end
          if ((st_res_2_15 == 3)) begin
            // clears sub states
            st_res_2_15 <= 0;
          end
          if ((st_res_2_15 == 3)) begin
          st_2 <= `S_2_121;
          end
        end
        `S_2_121: begin
          arg_15_389 <= r6_transform_264_338;
          st_2 <= `S_2_297;
        end
        `S_2_122: begin
          r4_transform_265_339 <= r1_bswap_16_397;
          st_2 <= `S_2_125;
        end
        `S_2_125: begin
          sram_addr_21 <= r0_transform_262_336;
          sram_wdata_21 <= r4_transform_265_339;
          st_2 <= `S_2_126;
        end
        `S_2_126: begin
          r0_transform_262_336 <= insn_o_2_166_0;
          st_2 <= `S_2_114;
        end
        `S_2_128: begin
          st_2 <= `S_2_129;
        end
        `S_2_129: begin
          r0_transform_262_336 <= 32'd16;
          st_2 <= `S_2_130;
        end
        `S_2_130: begin
          st_2 <= `S_2_131;
        end
        `S_2_131: begin
          r12_transform_266_340 <= insn_o_2_173_0;
          st_2 <= `S_2_132;
        end
        `S_2_132: begin
          if (r12_transform_266_340) begin
            st_2 <= `S_2_133;
          end else begin
            st_2 <= `S_2_167;
          end
        end
        `S_2_133: begin
          st_2 <= `S_2_135;
        end
        `S_2_135: begin
          r19_transform_267_341 <= insn_o_2_178_0;
          st_2 <= `S_2_138;
        end
        `S_2_138: begin
          sram_addr_21 <= r19_transform_267_341;
          st_2 <= `S_2_15;
        end
        `S_2_15: begin
          r21_transform_268_342 <= insn_o_2_66_0;
          st_2 <= `S_2_139;
        end
        `S_2_139: begin
          x_233_398 <= r21_transform_268_342;
          st_2 <= `S_2_317;
        end
        `S_2_140: begin
          r17_transform_269_343 <= r1_s1_234_404;
          st_2 <= `S_2_142;
        end
        `S_2_142: begin
          r24_transform_270_344 <= insn_o_2_190_0;
          st_2 <= `S_2_145;
        end
        `S_2_145: begin
          sram_addr_21 <= r24_transform_270_344;
          st_2 <= `S_2_16;
        end
        `S_2_16: begin
          r26_transform_271_345 <= insn_o_2_72_0;
          st_2 <= `S_2_146;
        end
        `S_2_146: begin
          r16_transform_272_346 <= insn_o_2_196_0;
          st_2 <= `S_2_149;
        end
        `S_2_149: begin
          r31_transform_273_347 <= insn_o_2_200_0;
          st_2 <= `S_2_152;
        end
        `S_2_152: begin
          sram_addr_21 <= r31_transform_273_347;
          st_2 <= `S_2_17;
        end
        `S_2_17: begin
          r33_transform_274_348 <= insn_o_2_75_0;
          st_2 <= `S_2_153;
        end
        `S_2_153: begin
          x_226_415 <= r33_transform_274_348;
          st_2 <= `S_2_359;
        end
        `S_2_154: begin
          r29_transform_275_349 <= r1_s0_227_421;
          st_2 <= `S_2_155;
        end
        `S_2_155: begin
          r15_transform_276_350 <= insn_o_2_211_0;
          st_2 <= `S_2_157;
        end
        `S_2_157: begin
          r36_transform_277_351 <= insn_o_2_214_0;
          st_2 <= `S_2_160;
        end
        `S_2_160: begin
          sram_addr_21 <= r36_transform_277_351;
          st_2 <= `S_2_18;
        end
        `S_2_18: begin
          r38_transform_278_352 <= insn_o_2_81_0;
          st_2 <= `S_2_161;
        end
        `S_2_161: begin
          r14_transform_279_353 <= insn_o_2_220_0;
          st_2 <= `S_2_164;
        end
        `S_2_164: begin
          sram_addr_21 <= r0_transform_262_336;
          sram_wdata_21 <= r14_transform_279_353;
          st_2 <= `S_2_165;
        end
        `S_2_165: begin
          r0_transform_262_336 <= insn_o_2_226_0;
          st_2 <= `S_2_130;
        end
        `S_2_167: begin
          st_2 <= `S_2_170;
        end
        `S_2_170: begin
          sram_addr_2 <= 32'd0;
          st_2 <= `S_2_22;
        end
        `S_2_22: begin
          r52_transform_280_354 <= insn_o_2_90_0;
          st_2 <= `S_2_171;
        end
        `S_2_171: begin
          r43_transform_281_355 <= r52_transform_280_354;
          st_2 <= `S_2_175;
        end
        `S_2_175: begin
          sram_addr_2 <= 32'd1;
          st_2 <= `S_2_24;
        end
        `S_2_24: begin
          r56_transform_282_356 <= insn_o_2_94_0;
          st_2 <= `S_2_176;
        end
        `S_2_176: begin
          r44_transform_283_357 <= r56_transform_282_356;
          st_2 <= `S_2_180;
        end
        `S_2_180: begin
          sram_addr_2 <= 32'd2;
          st_2 <= `S_2_25;
        end
        `S_2_25: begin
          r60_transform_284_358 <= insn_o_2_97_0;
          st_2 <= `S_2_181;
        end
        `S_2_181: begin
          r45_transform_285_359 <= r60_transform_284_358;
          st_2 <= `S_2_185;
        end
        `S_2_185: begin
          sram_addr_2 <= 32'd3;
          st_2 <= `S_2_27;
        end
        `S_2_27: begin
          r64_transform_286_360 <= insn_o_2_101_0;
          st_2 <= `S_2_186;
        end
        `S_2_186: begin
          r46_transform_287_361 <= r64_transform_286_360;
          st_2 <= `S_2_190;
        end
        `S_2_190: begin
          sram_addr_2 <= 32'd4;
          st_2 <= `S_2_28;
        end
        `S_2_28: begin
          r68_transform_288_362 <= insn_o_2_105_0;
          st_2 <= `S_2_191;
        end
        `S_2_191: begin
          r47_transform_289_363 <= r68_transform_288_362;
          st_2 <= `S_2_195;
        end
        `S_2_195: begin
          sram_addr_2 <= 32'd5;
          st_2 <= `S_2_29;
        end
        `S_2_29: begin
          r72_transform_290_364 <= insn_o_2_108_0;
          st_2 <= `S_2_196;
        end
        `S_2_196: begin
          r48_transform_291_365 <= r72_transform_290_364;
          st_2 <= `S_2_200;
        end
        `S_2_200: begin
          sram_addr_2 <= 32'd6;
          st_2 <= `S_2_32;
        end
        `S_2_32: begin
          r76_transform_292_366 <= insn_o_2_112_0;
          st_2 <= `S_2_201;
        end
        `S_2_201: begin
          r49_transform_293_367 <= r76_transform_292_366;
          st_2 <= `S_2_205;
        end
        `S_2_205: begin
          sram_addr_2 <= 32'd7;
          st_2 <= `S_2_33;
        end
        `S_2_33: begin
          r80_transform_294_368 <= insn_o_2_115_0;
          st_2 <= `S_2_206;
        end
        `S_2_206: begin
          r50_transform_295_369 <= r80_transform_294_368;
          st_2 <= `S_2_208;
        end
        `S_2_208: begin
          r0_transform_262_336 <= 32'd0;
          st_2 <= `S_2_209;
        end
        `S_2_209: begin
          st_2 <= `S_2_210;
        end
        `S_2_210: begin
          r84_transform_296_370 <= insn_o_2_289_0;
          st_2 <= `S_2_211;
        end
        `S_2_211: begin
          if (r84_transform_296_370) begin
            st_2 <= `S_2_212;
          end else begin
            st_2 <= `S_2_219;
          end
        end
        `S_2_212: begin
          st_2 <= `S_2_213;
        end
        `S_2_213: begin
          a_39_446 <= r43_transform_281_355;
          b_40_448 <= r44_transform_283_357;
          c_41_449 <= r45_transform_285_359;
          d_42_453 <= r46_transform_287_361;
          e_43_432 <= r47_transform_289_363;
          f_44_436 <= r48_transform_291_365;
          g_45_437 <= r49_transform_293_367;
          h_46_434 <= r50_transform_295_369;
          idx_47_440 <= r0_transform_262_336;
          st_2 <= `S_2_401;
        end
        `S_2_214: begin
          r43_transform_281_355 <= r9_iterate_48_561;
          r44_transform_283_357 <= r10_iterate_49_562;
          r45_transform_285_359 <= r11_iterate_50_563;
          r46_transform_287_361 <= r12_iterate_51_564;
          r47_transform_289_363 <= r13_iterate_52_565;
          r48_transform_291_365 <= r14_iterate_53_566;
          r49_transform_293_367 <= r15_iterate_54_567;
          r50_transform_295_369 <= r16_iterate_55_568;
          st_2 <= `S_2_216;
        end
        `S_2_216: begin
          r88_transform_297_371 <= insn_o_2_314_0;
          st_2 <= `S_2_217;
        end
        `S_2_217: begin
          r0_transform_262_336 <= r88_transform_297_371;
          st_2 <= `S_2_209;
        end
        `S_2_219: begin
          st_2 <= `S_2_222;
        end
        `S_2_222: begin
          sram_addr_2 <= 32'd0;
          st_2 <= `S_2_34;
        end
        `S_2_34: begin
          r90_transform_298_372 <= insn_o_2_119_0;
          st_2 <= `S_2_223;
        end
        `S_2_223: begin
          r93_transform_299_373 <= insn_o_2_324_0;
          st_2 <= `S_2_227;
        end
        `S_2_227: begin
          sram_addr_2 <= 32'd0;
          sram_wdata_2 <= r93_transform_299_373;
          st_2 <= `S_2_231;
        end
        `S_2_231: begin
          sram_addr_2 <= 32'd1;
          st_2 <= `S_2_37;
        end
        `S_2_37: begin
          r98_transform_300_374 <= insn_o_2_124_0;
          st_2 <= `S_2_232;
        end
        `S_2_232: begin
          r101_transform_301_375 <= insn_o_2_336_0;
          st_2 <= `S_2_236;
        end
        `S_2_236: begin
          sram_addr_2 <= 32'd1;
          sram_wdata_2 <= r101_transform_301_375;
          st_2 <= `S_2_240;
        end
        `S_2_240: begin
          sram_addr_2 <= 32'd2;
          st_2 <= `S_2_38;
        end
        `S_2_38: begin
          r106_transform_302_376 <= insn_o_2_129_0;
          st_2 <= `S_2_241;
        end
        `S_2_241: begin
          r109_transform_303_377 <= insn_o_2_348_0;
          st_2 <= `S_2_245;
        end
        `S_2_245: begin
          sram_addr_2 <= 32'd2;
          sram_wdata_2 <= r109_transform_303_377;
          st_2 <= `S_2_249;
        end
        `S_2_249: begin
          sram_addr_2 <= 32'd3;
          st_2 <= `S_2_39;
        end
        `S_2_39: begin
          r114_transform_304_378 <= insn_o_2_133_0;
          st_2 <= `S_2_250;
        end
        `S_2_250: begin
          r117_transform_305_379 <= insn_o_2_360_0;
          st_2 <= `S_2_254;
        end
        `S_2_254: begin
          sram_addr_2 <= 32'd3;
          sram_wdata_2 <= r117_transform_305_379;
          st_2 <= `S_2_258;
        end
        `S_2_258: begin
          sram_addr_2 <= 32'd4;
          st_2 <= `S_2_42;
        end
        `S_2_42: begin
          r122_transform_306_380 <= insn_o_2_138_0;
          st_2 <= `S_2_259;
        end
        `S_2_259: begin
          r125_transform_307_381 <= insn_o_2_372_0;
          st_2 <= `S_2_263;
        end
        `S_2_263: begin
          sram_addr_2 <= 32'd4;
          sram_wdata_2 <= r125_transform_307_381;
          st_2 <= `S_2_267;
        end
        `S_2_267: begin
          sram_addr_2 <= 32'd5;
          st_2 <= `S_2_43;
        end
        `S_2_43: begin
          r130_transform_308_382 <= insn_o_2_143_0;
          st_2 <= `S_2_268;
        end
        `S_2_268: begin
          r133_transform_309_383 <= insn_o_2_384_0;
          st_2 <= `S_2_272;
        end
        `S_2_272: begin
          sram_addr_2 <= 32'd5;
          sram_wdata_2 <= r133_transform_309_383;
          st_2 <= `S_2_276;
        end
        `S_2_276: begin
          sram_addr_2 <= 32'd6;
          st_2 <= `S_2_44;
        end
        `S_2_44: begin
          r138_transform_310_384 <= insn_o_2_154_0;
          st_2 <= `S_2_277;
        end
        `S_2_277: begin
          r141_transform_311_385 <= insn_o_2_396_0;
          st_2 <= `S_2_281;
        end
        `S_2_281: begin
          sram_addr_2 <= 32'd6;
          sram_wdata_2 <= r141_transform_311_385;
          st_2 <= `S_2_285;
        end
        `S_2_285: begin
          sram_addr_2 <= 32'd7;
          st_2 <= `S_2_47;
        end
        `S_2_47: begin
          r146_transform_312_386 <= insn_o_2_164_0;
          st_2 <= `S_2_286;
        end
        `S_2_286: begin
          r149_transform_313_387 <= insn_o_2_408_0;
          st_2 <= `S_2_290;
        end
        `S_2_290: begin
          sram_addr_2 <= 32'd7;
          sram_wdata_2 <= r149_transform_313_387;
          st_2 <= `S_2_19;
        end
        `S_2_297: begin
          r5_bswap_17_390 <= insn_o_2_421_0;
          st_2 <= `S_2_300;
        end
        `S_2_300: begin
          r8_bswap_18_391 <= insn_o_2_425_0;
          st_2 <= `S_2_301;
        end
        `S_2_301: begin
          r4_bswap_19_392 <= insn_o_2_427_0;
          st_2 <= `S_2_304;
        end
        `S_2_304: begin
          r11_bswap_20_393 <= insn_o_2_431_0;
          st_2 <= `S_2_305;
        end
        `S_2_305: begin
          r3_bswap_21_394 <= insn_o_2_433_0;
          st_2 <= `S_2_308;
        end
        `S_2_308: begin
          r14_bswap_22_395 <= insn_o_2_437_0;
          st_2 <= `S_2_309;
        end
        `S_2_309: begin
          r2_bswap_23_396 <= insn_o_2_439_0;
          st_2 <= `S_2_310;
        end
        `S_2_310: begin
          r1_bswap_16_397 <= r2_bswap_23_396;
          st_2 <= `S_2_122;
        end
        `S_2_317: begin
          arg_186_405 <= x_233_398;
          st_2 <= `S_2_334;
        end
        `S_2_318: begin
          r4_s1_235_399 <= r1_ror32_17_187_409;
          st_2 <= `S_2_320;
        end
        `S_2_320: begin
          arg_196_410 <= x_233_398;
          st_2 <= `S_2_347;
        end
        `S_2_321: begin
          r6_s1_236_400 <= r1_ror32_19_197_414;
          st_2 <= `S_2_322;
        end
        `S_2_322: begin
          r3_s1_237_401 <= insn_o_2_460_0;
          st_2 <= `S_2_324;
        end
        `S_2_324: begin
          r8_s1_238_402 <= insn_o_2_463_0;
          st_2 <= `S_2_325;
        end
        `S_2_325: begin
          r2_s1_239_403 <= insn_o_2_465_0;
          st_2 <= `S_2_326;
        end
        `S_2_326: begin
          r1_s1_234_404 <= r2_s1_239_403;
          st_2 <= `S_2_140;
        end
        `S_2_334: begin
          r3_ror32_17_188_406 <= insn_o_2_476_0;
          st_2 <= `S_2_337;
        end
        `S_2_337: begin
          r6_ror32_17_189_407 <= insn_o_2_480_0;
          st_2 <= `S_2_338;
        end
        `S_2_338: begin
          r2_ror32_17_190_408 <= insn_o_2_482_0;
          st_2 <= `S_2_339;
        end
        `S_2_339: begin
          r1_ror32_17_187_409 <= r2_ror32_17_190_408;
          st_2 <= `S_2_318;
        end
        `S_2_347: begin
          r3_ror32_19_198_411 <= insn_o_2_493_0;
          st_2 <= `S_2_350;
        end
        `S_2_350: begin
          r6_ror32_19_199_412 <= insn_o_2_497_0;
          st_2 <= `S_2_351;
        end
        `S_2_351: begin
          r2_ror32_19_200_413 <= insn_o_2_499_0;
          st_2 <= `S_2_352;
        end
        `S_2_352: begin
          r1_ror32_19_197_414 <= r2_ror32_19_200_413;
          st_2 <= `S_2_321;
        end
        `S_2_359: begin
          arg_221_422 <= x_226_415;
          st_2 <= `S_2_376;
        end
        `S_2_360: begin
          r4_s0_228_416 <= r1_ror32_7_222_426;
          st_2 <= `S_2_362;
        end
        `S_2_362: begin
          arg_191_427 <= x_226_415;
          st_2 <= `S_2_389;
        end
        `S_2_363: begin
          r6_s0_229_417 <= r1_ror32_18_192_431;
          st_2 <= `S_2_364;
        end
        `S_2_364: begin
          r3_s0_230_418 <= insn_o_2_520_0;
          st_2 <= `S_2_366;
        end
        `S_2_366: begin
          r8_s0_231_419 <= insn_o_2_523_0;
          st_2 <= `S_2_367;
        end
        `S_2_367: begin
          r2_s0_232_420 <= insn_o_2_525_0;
          st_2 <= `S_2_368;
        end
        `S_2_368: begin
          r1_s0_227_421 <= r2_s0_232_420;
          st_2 <= `S_2_154;
        end
        `S_2_376: begin
          r3_ror32_7_223_423 <= insn_o_2_536_0;
          st_2 <= `S_2_379;
        end
        `S_2_379: begin
          r6_ror32_7_224_424 <= insn_o_2_540_0;
          st_2 <= `S_2_380;
        end
        `S_2_380: begin
          r2_ror32_7_225_425 <= insn_o_2_542_0;
          st_2 <= `S_2_381;
        end
        `S_2_381: begin
          r1_ror32_7_222_426 <= r2_ror32_7_225_425;
          st_2 <= `S_2_360;
        end
        `S_2_389: begin
          r3_ror32_18_193_428 <= insn_o_2_553_0;
          st_2 <= `S_2_392;
        end
        `S_2_392: begin
          r6_ror32_18_194_429 <= insn_o_2_557_0;
          st_2 <= `S_2_393;
        end
        `S_2_393: begin
          r2_ror32_18_195_430 <= insn_o_2_559_0;
          st_2 <= `S_2_394;
        end
        `S_2_394: begin
          r1_ror32_18_192_431 <= r2_ror32_18_195_430;
          st_2 <= `S_2_363;
        end
        `S_2_401: begin
          x_31_569 <= e_43_432;
          st_2 <= `S_2_674;
        end
        `S_2_402: begin
          r23_iterate_56_433 <= r1_e1_32_575;
          st_2 <= `S_2_403;
        end
        `S_2_403: begin
          r22_iterate_57_435 <= insn_o_2_574_0;
          st_2 <= `S_2_405;
        end
        `S_2_405: begin
          x_0_594 <= e_43_432;
          y_1_591 <= f_44_436;
          z_2_592 <= g_45_437;
          st_2 <= `S_2_729;
        end
        `S_2_406: begin
          r25_iterate_58_438 <= r3_Ch_3_597;
          st_2 <= `S_2_407;
        end
        `S_2_407: begin
          r21_iterate_59_439 <= insn_o_2_584_0;
          st_2 <= `S_2_410;
        end
        `S_2_410: begin
          sram_addr_20 <= idx_47_440;
          st_2 <= `S_2_48;
        end
        `S_2_48: begin
          r27_iterate_60_441 <= insn_o_2_181_0;
          st_2 <= `S_2_411;
        end
        `S_2_411: begin
          r20_iterate_61_442 <= insn_o_2_590_0;
          st_2 <= `S_2_414;
        end
        `S_2_414: begin
          sram_addr_21 <= idx_47_440;
          st_2 <= `S_2_49;
        end
        `S_2_49: begin
          r30_iterate_62_443 <= insn_o_2_189_0;
          st_2 <= `S_2_415;
        end
        `S_2_415: begin
          r19_iterate_63_444 <= insn_o_2_596_0;
          st_2 <= `S_2_416;
        end
        `S_2_416: begin
          r17_iterate_64_445 <= r19_iterate_63_444;
          st_2 <= `S_2_418;
        end
        `S_2_418: begin
          x_24_598 <= a_39_446;
          st_2 <= `S_2_739;
        end
        `S_2_419: begin
          r34_iterate_65_447 <= r1_e0_25_604;
          st_2 <= `S_2_421;
        end
        `S_2_421: begin
          x_7_620 <= a_39_446;
          y_8_621 <= b_40_448;
          z_9_624 <= c_41_449;
          st_2 <= `S_2_794;
        end
        `S_2_422: begin
          r36_iterate_66_450 <= r3_Maj_10_627;
          st_2 <= `S_2_423;
        end
        `S_2_423: begin
          r33_iterate_67_451 <= insn_o_2_614_0;
          st_2 <= `S_2_424;
        end
        `S_2_424: begin
          r18_iterate_68_452 <= r33_iterate_67_451;
          st_2 <= `S_2_425;
        end
        `S_2_425: begin
          r38_iterate_69_454 <= insn_o_2_618_0;
          st_2 <= `S_2_426;
        end
        `S_2_426: begin
          d_42_453 <= r38_iterate_69_454;
          st_2 <= `S_2_427;
        end
        `S_2_427: begin
          r39_iterate_70_455 <= insn_o_2_622_0;
          st_2 <= `S_2_428;
        end
        `S_2_428: begin
          h_46_434 <= r39_iterate_70_455;
          st_2 <= `S_2_430;
        end
        `S_2_430: begin
          x_31_628 <= d_42_453;
          st_2 <= `S_2_805;
        end
        `S_2_431: begin
          r44_iterate_71_456 <= r1_e1_32_634;
          st_2 <= `S_2_432;
        end
        `S_2_432: begin
          r43_iterate_72_457 <= insn_o_2_632_0;
          st_2 <= `S_2_434;
        end
        `S_2_434: begin
          x_0_653 <= d_42_453;
          y_1_650 <= e_43_432;
          z_2_651 <= f_44_436;
          st_2 <= `S_2_860;
        end
        `S_2_435: begin
          r46_iterate_73_458 <= r3_Ch_3_656;
          st_2 <= `S_2_436;
        end
        `S_2_436: begin
          r42_iterate_74_459 <= insn_o_2_642_0;
          st_2 <= `S_2_438;
        end
        `S_2_438: begin
          r48_iterate_75_460 <= insn_o_2_645_0;
          st_2 <= `S_2_441;
        end
        `S_2_441: begin
          sram_addr_20 <= r48_iterate_75_460;
          st_2 <= `S_2_52;
        end
        `S_2_52: begin
          r50_iterate_76_461 <= insn_o_2_194_0;
          st_2 <= `S_2_442;
        end
        `S_2_442: begin
          r41_iterate_77_462 <= insn_o_2_651_0;
          st_2 <= `S_2_444;
        end
        `S_2_444: begin
          r53_iterate_78_463 <= insn_o_2_654_0;
          st_2 <= `S_2_447;
        end
        `S_2_447: begin
          sram_addr_21 <= r53_iterate_78_463;
          st_2 <= `S_2_53;
        end
        `S_2_53: begin
          r55_iterate_79_464 <= insn_o_2_202_0;
          st_2 <= `S_2_448;
        end
        `S_2_448: begin
          r40_iterate_80_465 <= insn_o_2_660_0;
          st_2 <= `S_2_449;
        end
        `S_2_449: begin
          r17_iterate_64_445 <= r40_iterate_80_465;
          st_2 <= `S_2_451;
        end
        `S_2_451: begin
          x_24_657 <= h_46_434;
          st_2 <= `S_2_870;
        end
        `S_2_452: begin
          r59_iterate_81_466 <= r1_e0_25_663;
          st_2 <= `S_2_454;
        end
        `S_2_454: begin
          x_7_679 <= h_46_434;
          y_8_680 <= a_39_446;
          z_9_683 <= b_40_448;
          st_2 <= `S_2_925;
        end
        `S_2_455: begin
          r61_iterate_82_467 <= r3_Maj_10_686;
          st_2 <= `S_2_456;
        end
        `S_2_456: begin
          r58_iterate_83_468 <= insn_o_2_678_0;
          st_2 <= `S_2_457;
        end
        `S_2_457: begin
          r18_iterate_68_452 <= r58_iterate_83_468;
          st_2 <= `S_2_458;
        end
        `S_2_458: begin
          r63_iterate_84_469 <= insn_o_2_682_0;
          st_2 <= `S_2_459;
        end
        `S_2_459: begin
          c_41_449 <= r63_iterate_84_469;
          st_2 <= `S_2_460;
        end
        `S_2_460: begin
          r64_iterate_85_470 <= insn_o_2_686_0;
          st_2 <= `S_2_461;
        end
        `S_2_461: begin
          g_45_437 <= r64_iterate_85_470;
          st_2 <= `S_2_463;
        end
        `S_2_463: begin
          x_31_687 <= c_41_449;
          st_2 <= `S_2_936;
        end
        `S_2_464: begin
          r69_iterate_86_471 <= r1_e1_32_693;
          st_2 <= `S_2_465;
        end
        `S_2_465: begin
          r68_iterate_87_472 <= insn_o_2_696_0;
          st_2 <= `S_2_467;
        end
        `S_2_467: begin
          x_0_712 <= c_41_449;
          y_1_709 <= d_42_453;
          z_2_710 <= e_43_432;
          st_2 <= `S_2_991;
        end
        `S_2_468: begin
          r71_iterate_88_473 <= r3_Ch_3_715;
          st_2 <= `S_2_469;
        end
        `S_2_469: begin
          r67_iterate_89_474 <= insn_o_2_706_0;
          st_2 <= `S_2_471;
        end
        `S_2_471: begin
          r73_iterate_90_475 <= insn_o_2_709_0;
          st_2 <= `S_2_474;
        end
        `S_2_474: begin
          sram_addr_20 <= r73_iterate_90_475;
          st_2 <= `S_2_54;
        end
        `S_2_54: begin
          r75_iterate_91_476 <= insn_o_2_206_0;
          st_2 <= `S_2_475;
        end
        `S_2_475: begin
          r66_iterate_92_477 <= insn_o_2_715_0;
          st_2 <= `S_2_477;
        end
        `S_2_477: begin
          r78_iterate_93_478 <= insn_o_2_718_0;
          st_2 <= `S_2_480;
        end
        `S_2_480: begin
          sram_addr_21 <= r78_iterate_93_478;
          st_2 <= `S_2_57;
        end
        `S_2_57: begin
          r80_iterate_94_479 <= insn_o_2_217_0;
          st_2 <= `S_2_481;
        end
        `S_2_481: begin
          r65_iterate_95_480 <= insn_o_2_724_0;
          st_2 <= `S_2_482;
        end
        `S_2_482: begin
          r17_iterate_64_445 <= r65_iterate_95_480;
          st_2 <= `S_2_484;
        end
        `S_2_484: begin
          x_24_716 <= g_45_437;
          st_2 <= `S_2_1001;
        end
        `S_2_485: begin
          r84_iterate_96_481 <= r1_e0_25_722;
          st_2 <= `S_2_487;
        end
        `S_2_487: begin
          x_7_738 <= g_45_437;
          y_8_739 <= h_46_434;
          z_9_742 <= a_39_446;
          st_2 <= `S_2_1056;
        end
        `S_2_488: begin
          r86_iterate_97_482 <= r3_Maj_10_745;
          st_2 <= `S_2_489;
        end
        `S_2_489: begin
          r83_iterate_98_483 <= insn_o_2_742_0;
          st_2 <= `S_2_490;
        end
        `S_2_490: begin
          r18_iterate_68_452 <= r83_iterate_98_483;
          st_2 <= `S_2_491;
        end
        `S_2_491: begin
          r88_iterate_99_484 <= insn_o_2_746_0;
          st_2 <= `S_2_492;
        end
        `S_2_492: begin
          b_40_448 <= r88_iterate_99_484;
          st_2 <= `S_2_493;
        end
        `S_2_493: begin
          r89_iterate_100_485 <= insn_o_2_750_0;
          st_2 <= `S_2_494;
        end
        `S_2_494: begin
          f_44_436 <= r89_iterate_100_485;
          st_2 <= `S_2_496;
        end
        `S_2_496: begin
          x_31_746 <= b_40_448;
          st_2 <= `S_2_1067;
        end
        `S_2_497: begin
          r94_iterate_101_486 <= r1_e1_32_752;
          st_2 <= `S_2_498;
        end
        `S_2_498: begin
          r93_iterate_102_487 <= insn_o_2_760_0;
          st_2 <= `S_2_500;
        end
        `S_2_500: begin
          x_0_771 <= b_40_448;
          y_1_768 <= c_41_449;
          z_2_769 <= d_42_453;
          st_2 <= `S_2_1122;
        end
        `S_2_501: begin
          r96_iterate_103_488 <= r3_Ch_3_774;
          st_2 <= `S_2_502;
        end
        `S_2_502: begin
          r92_iterate_104_489 <= insn_o_2_770_0;
          st_2 <= `S_2_504;
        end
        `S_2_504: begin
          r98_iterate_105_490 <= insn_o_2_773_0;
          st_2 <= `S_2_507;
        end
        `S_2_507: begin
          sram_addr_20 <= r98_iterate_105_490;
          st_2 <= `S_2_58;
        end
        `S_2_58: begin
          r100_iterate_106_491 <= insn_o_2_223_0;
          st_2 <= `S_2_508;
        end
        `S_2_508: begin
          r91_iterate_107_492 <= insn_o_2_779_0;
          st_2 <= `S_2_510;
        end
        `S_2_510: begin
          r103_iterate_108_493 <= insn_o_2_782_0;
          st_2 <= `S_2_513;
        end
        `S_2_513: begin
          sram_addr_21 <= r103_iterate_108_493;
          st_2 <= `S_2_59;
        end
        `S_2_59: begin
          r105_iterate_109_494 <= insn_o_2_230_0;
          st_2 <= `S_2_514;
        end
        `S_2_514: begin
          r90_iterate_110_495 <= insn_o_2_788_0;
          st_2 <= `S_2_515;
        end
        `S_2_515: begin
          r17_iterate_64_445 <= r90_iterate_110_495;
          st_2 <= `S_2_517;
        end
        `S_2_517: begin
          x_24_775 <= f_44_436;
          st_2 <= `S_2_1132;
        end
        `S_2_518: begin
          r109_iterate_111_496 <= r1_e0_25_781;
          st_2 <= `S_2_520;
        end
        `S_2_520: begin
          x_7_797 <= f_44_436;
          y_8_798 <= g_45_437;
          z_9_801 <= h_46_434;
          st_2 <= `S_2_1187;
        end
        `S_2_521: begin
          r111_iterate_112_497 <= r3_Maj_10_804;
          st_2 <= `S_2_522;
        end
        `S_2_522: begin
          r108_iterate_113_498 <= insn_o_2_806_0;
          st_2 <= `S_2_523;
        end
        `S_2_523: begin
          r18_iterate_68_452 <= r108_iterate_113_498;
          st_2 <= `S_2_524;
        end
        `S_2_524: begin
          r113_iterate_114_499 <= insn_o_2_810_0;
          st_2 <= `S_2_525;
        end
        `S_2_525: begin
          a_39_446 <= r113_iterate_114_499;
          st_2 <= `S_2_526;
        end
        `S_2_526: begin
          r114_iterate_115_500 <= insn_o_2_814_0;
          st_2 <= `S_2_527;
        end
        `S_2_527: begin
          e_43_432 <= r114_iterate_115_500;
          st_2 <= `S_2_529;
        end
        `S_2_529: begin
          x_31_805 <= a_39_446;
          st_2 <= `S_2_1198;
        end
        `S_2_530: begin
          r119_iterate_116_501 <= r1_e1_32_811;
          st_2 <= `S_2_531;
        end
        `S_2_531: begin
          r118_iterate_117_502 <= insn_o_2_824_0;
          st_2 <= `S_2_533;
        end
        `S_2_533: begin
          x_0_830 <= a_39_446;
          y_1_827 <= b_40_448;
          z_2_828 <= c_41_449;
          st_2 <= `S_2_1253;
        end
        `S_2_534: begin
          r121_iterate_118_503 <= r3_Ch_3_833;
          st_2 <= `S_2_535;
        end
        `S_2_535: begin
          r117_iterate_119_504 <= insn_o_2_834_0;
          st_2 <= `S_2_537;
        end
        `S_2_537: begin
          r123_iterate_120_505 <= insn_o_2_837_0;
          st_2 <= `S_2_540;
        end
        `S_2_540: begin
          sram_addr_20 <= r123_iterate_120_505;
          st_2 <= `S_2_63;
        end
        `S_2_63: begin
          r125_iterate_121_506 <= insn_o_2_236_0;
          st_2 <= `S_2_541;
        end
        `S_2_541: begin
          r116_iterate_122_507 <= insn_o_2_843_0;
          st_2 <= `S_2_543;
        end
        `S_2_543: begin
          r128_iterate_123_508 <= insn_o_2_846_0;
          st_2 <= `S_2_546;
        end
        `S_2_546: begin
          sram_addr_21 <= r128_iterate_123_508;
          st_2 <= `S_2_64;
        end
        `S_2_64: begin
          r130_iterate_124_509 <= insn_o_2_239_0;
          st_2 <= `S_2_547;
        end
        `S_2_547: begin
          r115_iterate_125_510 <= insn_o_2_852_0;
          st_2 <= `S_2_548;
        end
        `S_2_548: begin
          r17_iterate_64_445 <= r115_iterate_125_510;
          st_2 <= `S_2_550;
        end
        `S_2_550: begin
          x_24_834 <= e_43_432;
          st_2 <= `S_2_1263;
        end
        `S_2_551: begin
          r134_iterate_126_511 <= r1_e0_25_840;
          st_2 <= `S_2_553;
        end
        `S_2_553: begin
          x_7_856 <= e_43_432;
          y_8_857 <= f_44_436;
          z_9_860 <= g_45_437;
          st_2 <= `S_2_1318;
        end
        `S_2_554: begin
          r136_iterate_127_512 <= r3_Maj_10_863;
          st_2 <= `S_2_555;
        end
        `S_2_555: begin
          r133_iterate_128_513 <= insn_o_2_870_0;
          st_2 <= `S_2_556;
        end
        `S_2_556: begin
          r18_iterate_68_452 <= r133_iterate_128_513;
          st_2 <= `S_2_557;
        end
        `S_2_557: begin
          r138_iterate_129_514 <= insn_o_2_874_0;
          st_2 <= `S_2_558;
        end
        `S_2_558: begin
          h_46_434 <= r138_iterate_129_514;
          st_2 <= `S_2_559;
        end
        `S_2_559: begin
          r139_iterate_130_515 <= insn_o_2_878_0;
          st_2 <= `S_2_560;
        end
        `S_2_560: begin
          d_42_453 <= r139_iterate_130_515;
          st_2 <= `S_2_562;
        end
        `S_2_562: begin
          x_31_864 <= h_46_434;
          st_2 <= `S_2_1329;
        end
        `S_2_563: begin
          r144_iterate_131_516 <= r1_e1_32_870;
          st_2 <= `S_2_564;
        end
        `S_2_564: begin
          r143_iterate_132_517 <= insn_o_2_888_0;
          st_2 <= `S_2_566;
        end
        `S_2_566: begin
          x_0_889 <= h_46_434;
          y_1_886 <= a_39_446;
          z_2_887 <= b_40_448;
          st_2 <= `S_2_1384;
        end
        `S_2_567: begin
          r146_iterate_133_518 <= r3_Ch_3_892;
          st_2 <= `S_2_568;
        end
        `S_2_568: begin
          r142_iterate_134_519 <= insn_o_2_898_0;
          st_2 <= `S_2_570;
        end
        `S_2_570: begin
          r148_iterate_135_520 <= insn_o_2_901_0;
          st_2 <= `S_2_573;
        end
        `S_2_573: begin
          sram_addr_20 <= r148_iterate_135_520;
          st_2 <= `S_2_65;
        end
        `S_2_65: begin
          r150_iterate_136_521 <= insn_o_2_245_0;
          st_2 <= `S_2_574;
        end
        `S_2_574: begin
          r141_iterate_137_522 <= insn_o_2_907_0;
          st_2 <= `S_2_576;
        end
        `S_2_576: begin
          r153_iterate_138_523 <= insn_o_2_910_0;
          st_2 <= `S_2_579;
        end
        `S_2_579: begin
          sram_addr_21 <= r153_iterate_138_523;
          st_2 <= `S_2_67;
        end
        `S_2_67: begin
          r155_iterate_139_524 <= insn_o_2_251_0;
          st_2 <= `S_2_580;
        end
        `S_2_580: begin
          r140_iterate_140_525 <= insn_o_2_916_0;
          st_2 <= `S_2_581;
        end
        `S_2_581: begin
          r17_iterate_64_445 <= r140_iterate_140_525;
          st_2 <= `S_2_583;
        end
        `S_2_583: begin
          x_24_893 <= d_42_453;
          st_2 <= `S_2_1394;
        end
        `S_2_584: begin
          r159_iterate_141_526 <= r1_e0_25_899;
          st_2 <= `S_2_586;
        end
        `S_2_586: begin
          x_7_915 <= d_42_453;
          y_8_916 <= e_43_432;
          z_9_919 <= f_44_436;
          st_2 <= `S_2_1449;
        end
        `S_2_587: begin
          r161_iterate_142_527 <= r3_Maj_10_922;
          st_2 <= `S_2_588;
        end
        `S_2_588: begin
          r158_iterate_143_528 <= insn_o_2_934_0;
          st_2 <= `S_2_589;
        end
        `S_2_589: begin
          r18_iterate_68_452 <= r158_iterate_143_528;
          st_2 <= `S_2_590;
        end
        `S_2_590: begin
          r163_iterate_144_529 <= insn_o_2_938_0;
          st_2 <= `S_2_591;
        end
        `S_2_591: begin
          g_45_437 <= r163_iterate_144_529;
          st_2 <= `S_2_592;
        end
        `S_2_592: begin
          r164_iterate_145_530 <= insn_o_2_942_0;
          st_2 <= `S_2_593;
        end
        `S_2_593: begin
          c_41_449 <= r164_iterate_145_530;
          st_2 <= `S_2_595;
        end
        `S_2_595: begin
          x_31_923 <= g_45_437;
          st_2 <= `S_2_1460;
        end
        `S_2_596: begin
          r169_iterate_146_531 <= r1_e1_32_929;
          st_2 <= `S_2_597;
        end
        `S_2_597: begin
          r168_iterate_147_532 <= insn_o_2_952_0;
          st_2 <= `S_2_599;
        end
        `S_2_599: begin
          x_0_948 <= g_45_437;
          y_1_945 <= h_46_434;
          z_2_946 <= a_39_446;
          st_2 <= `S_2_1515;
        end
        `S_2_600: begin
          r171_iterate_148_533 <= r3_Ch_3_951;
          st_2 <= `S_2_601;
        end
        `S_2_601: begin
          r167_iterate_149_534 <= insn_o_2_962_0;
          st_2 <= `S_2_603;
        end
        `S_2_603: begin
          r173_iterate_150_535 <= insn_o_2_965_0;
          st_2 <= `S_2_606;
        end
        `S_2_606: begin
          sram_addr_20 <= r173_iterate_150_535;
          st_2 <= `S_2_68;
        end
        `S_2_68: begin
          r175_iterate_151_536 <= insn_o_2_257_0;
          st_2 <= `S_2_607;
        end
        `S_2_607: begin
          r166_iterate_152_537 <= insn_o_2_971_0;
          st_2 <= `S_2_609;
        end
        `S_2_609: begin
          r178_iterate_153_538 <= insn_o_2_974_0;
          st_2 <= `S_2_612;
        end
        `S_2_612: begin
          sram_addr_21 <= r178_iterate_153_538;
          st_2 <= `S_2_69;
        end
        `S_2_69: begin
          r180_iterate_154_539 <= insn_o_2_260_0;
          st_2 <= `S_2_613;
        end
        `S_2_613: begin
          r165_iterate_155_540 <= insn_o_2_980_0;
          st_2 <= `S_2_614;
        end
        `S_2_614: begin
          r17_iterate_64_445 <= r165_iterate_155_540;
          st_2 <= `S_2_616;
        end
        `S_2_616: begin
          x_24_952 <= c_41_449;
          st_2 <= `S_2_1525;
        end
        `S_2_617: begin
          r184_iterate_156_541 <= r1_e0_25_958;
          st_2 <= `S_2_619;
        end
        `S_2_619: begin
          x_7_974 <= c_41_449;
          y_8_975 <= d_42_453;
          z_9_978 <= e_43_432;
          st_2 <= `S_2_1580;
        end
        `S_2_620: begin
          r186_iterate_157_542 <= r3_Maj_10_981;
          st_2 <= `S_2_621;
        end
        `S_2_621: begin
          r183_iterate_158_543 <= insn_o_2_998_0;
          st_2 <= `S_2_622;
        end
        `S_2_622: begin
          r18_iterate_68_452 <= r183_iterate_158_543;
          st_2 <= `S_2_623;
        end
        `S_2_623: begin
          r188_iterate_159_544 <= insn_o_2_1002_0;
          st_2 <= `S_2_624;
        end
        `S_2_624: begin
          f_44_436 <= r188_iterate_159_544;
          st_2 <= `S_2_625;
        end
        `S_2_625: begin
          r189_iterate_160_545 <= insn_o_2_1006_0;
          st_2 <= `S_2_626;
        end
        `S_2_626: begin
          b_40_448 <= r189_iterate_160_545;
          st_2 <= `S_2_628;
        end
        `S_2_628: begin
          x_31_982 <= f_44_436;
          st_2 <= `S_2_1591;
        end
        `S_2_629: begin
          r194_iterate_161_546 <= r1_e1_32_988;
          st_2 <= `S_2_630;
        end
        `S_2_630: begin
          r193_iterate_162_547 <= insn_o_2_1016_0;
          st_2 <= `S_2_632;
        end
        `S_2_632: begin
          x_0_1007 <= f_44_436;
          y_1_1004 <= g_45_437;
          z_2_1005 <= h_46_434;
          st_2 <= `S_2_1646;
        end
        `S_2_633: begin
          r196_iterate_163_548 <= r3_Ch_3_1010;
          st_2 <= `S_2_634;
        end
        `S_2_634: begin
          r192_iterate_164_549 <= insn_o_2_1026_0;
          st_2 <= `S_2_636;
        end
        `S_2_636: begin
          r198_iterate_165_550 <= insn_o_2_1029_0;
          st_2 <= `S_2_639;
        end
        `S_2_639: begin
          sram_addr_20 <= r198_iterate_165_550;
          st_2 <= `S_2_70;
        end
        `S_2_70: begin
          r200_iterate_166_551 <= insn_o_2_266_0;
          st_2 <= `S_2_640;
        end
        `S_2_640: begin
          r191_iterate_167_552 <= insn_o_2_1035_0;
          st_2 <= `S_2_642;
        end
        `S_2_642: begin
          r203_iterate_168_553 <= insn_o_2_1038_0;
          st_2 <= `S_2_645;
        end
        `S_2_645: begin
          sram_addr_21 <= r203_iterate_168_553;
          st_2 <= `S_2_71;
        end
        `S_2_71: begin
          r205_iterate_169_554 <= insn_o_2_272_0;
          st_2 <= `S_2_646;
        end
        `S_2_646: begin
          r190_iterate_170_555 <= insn_o_2_1044_0;
          st_2 <= `S_2_647;
        end
        `S_2_647: begin
          r17_iterate_64_445 <= r190_iterate_170_555;
          st_2 <= `S_2_649;
        end
        `S_2_649: begin
          x_24_1011 <= b_40_448;
          st_2 <= `S_2_1656;
        end
        `S_2_650: begin
          r209_iterate_171_556 <= r1_e0_25_1017;
          st_2 <= `S_2_652;
        end
        `S_2_652: begin
          x_7_1033 <= b_40_448;
          y_8_1034 <= c_41_449;
          z_9_1037 <= d_42_453;
          st_2 <= `S_2_1711;
        end
        `S_2_653: begin
          r211_iterate_172_557 <= r3_Maj_10_1040;
          st_2 <= `S_2_654;
        end
        `S_2_654: begin
          r208_iterate_173_558 <= insn_o_2_1062_0;
          st_2 <= `S_2_655;
        end
        `S_2_655: begin
          r18_iterate_68_452 <= r208_iterate_173_558;
          st_2 <= `S_2_656;
        end
        `S_2_656: begin
          r213_iterate_174_559 <= insn_o_2_1066_0;
          st_2 <= `S_2_657;
        end
        `S_2_657: begin
          e_43_432 <= r213_iterate_174_559;
          st_2 <= `S_2_658;
        end
        `S_2_658: begin
          r214_iterate_175_560 <= insn_o_2_1070_0;
          st_2 <= `S_2_659;
        end
        `S_2_659: begin
          a_39_446 <= r214_iterate_175_560;
          st_2 <= `S_2_660;
        end
        `S_2_660: begin
          r9_iterate_48_561 <= a_39_446;
          st_2 <= `S_2_661;
        end
        `S_2_661: begin
          r10_iterate_49_562 <= b_40_448;
          st_2 <= `S_2_662;
        end
        `S_2_662: begin
          r11_iterate_50_563 <= c_41_449;
          st_2 <= `S_2_663;
        end
        `S_2_663: begin
          r12_iterate_51_564 <= d_42_453;
          st_2 <= `S_2_664;
        end
        `S_2_664: begin
          r13_iterate_52_565 <= e_43_432;
          st_2 <= `S_2_665;
        end
        `S_2_665: begin
          r14_iterate_53_566 <= f_44_436;
          st_2 <= `S_2_666;
        end
        `S_2_666: begin
          r15_iterate_54_567 <= g_45_437;
          st_2 <= `S_2_667;
        end
        `S_2_667: begin
          r16_iterate_55_568 <= h_46_434;
          st_2 <= `S_2_214;
        end
        `S_2_674: begin
          arg_216_576 <= x_31_569;
          st_2 <= `S_2_692;
        end
        `S_2_675: begin
          r4_e1_33_570 <= r1_ror32_6_217_580;
          st_2 <= `S_2_677;
        end
        `S_2_677: begin
          arg_176_581 <= x_31_569;
          st_2 <= `S_2_705;
        end
        `S_2_678: begin
          r6_e1_34_571 <= r1_ror32_11_177_585;
          st_2 <= `S_2_679;
        end
        `S_2_679: begin
          r3_e1_35_572 <= insn_o_2_1107_0;
          st_2 <= `S_2_681;
        end
        `S_2_681: begin
          arg_211_586 <= x_31_569;
          st_2 <= `S_2_718;
        end
        `S_2_682: begin
          r8_e1_36_573 <= r1_ror32_25_212_590;
          st_2 <= `S_2_683;
        end
        `S_2_683: begin
          r2_e1_37_574 <= insn_o_2_1115_0;
          st_2 <= `S_2_684;
        end
        `S_2_684: begin
          r1_e1_32_575 <= r2_e1_37_574;
          st_2 <= `S_2_402;
        end
        `S_2_692: begin
          r3_ror32_6_218_577 <= insn_o_2_1126_0;
          st_2 <= `S_2_695;
        end
        `S_2_695: begin
          r6_ror32_6_219_578 <= insn_o_2_1130_0;
          st_2 <= `S_2_696;
        end
        `S_2_696: begin
          r2_ror32_6_220_579 <= insn_o_2_1132_0;
          st_2 <= `S_2_697;
        end
        `S_2_697: begin
          r1_ror32_6_217_580 <= r2_ror32_6_220_579;
          st_2 <= `S_2_675;
        end
        `S_2_705: begin
          r3_ror32_11_178_582 <= insn_o_2_1143_0;
          st_2 <= `S_2_708;
        end
        `S_2_708: begin
          r6_ror32_11_179_583 <= insn_o_2_1147_0;
          st_2 <= `S_2_709;
        end
        `S_2_709: begin
          r2_ror32_11_180_584 <= insn_o_2_1149_0;
          st_2 <= `S_2_710;
        end
        `S_2_710: begin
          r1_ror32_11_177_585 <= r2_ror32_11_180_584;
          st_2 <= `S_2_678;
        end
        `S_2_718: begin
          r3_ror32_25_213_587 <= insn_o_2_1160_0;
          st_2 <= `S_2_721;
        end
        `S_2_721: begin
          r6_ror32_25_214_588 <= insn_o_2_1164_0;
          st_2 <= `S_2_722;
        end
        `S_2_722: begin
          r2_ror32_25_215_589 <= insn_o_2_1166_0;
          st_2 <= `S_2_723;
        end
        `S_2_723: begin
          r1_ror32_25_212_590 <= r2_ror32_25_215_589;
          st_2 <= `S_2_682;
        end
        `S_2_729: begin
          r6_Ch_4_593 <= insn_o_2_1175_0;
          st_2 <= `S_2_730;
        end
        `S_2_730: begin
          r5_Ch_5_595 <= insn_o_2_1177_0;
          st_2 <= `S_2_731;
        end
        `S_2_731: begin
          r4_Ch_6_596 <= insn_o_2_1179_0;
          st_2 <= `S_2_732;
        end
        `S_2_732: begin
          r3_Ch_3_597 <= r4_Ch_6_596;
          st_2 <= `S_2_406;
        end
        `S_2_739: begin
          arg_201_605 <= x_24_598;
          st_2 <= `S_2_757;
        end
        `S_2_740: begin
          r4_e0_26_599 <= r1_ror32_2_202_609;
          st_2 <= `S_2_742;
        end
        `S_2_742: begin
          arg_181_610 <= x_24_598;
          st_2 <= `S_2_770;
        end
        `S_2_743: begin
          r6_e0_27_600 <= r1_ror32_13_182_614;
          st_2 <= `S_2_744;
        end
        `S_2_744: begin
          r3_e0_28_601 <= insn_o_2_1200_0;
          st_2 <= `S_2_746;
        end
        `S_2_746: begin
          arg_206_615 <= x_24_598;
          st_2 <= `S_2_783;
        end
        `S_2_747: begin
          r8_e0_29_602 <= r1_ror32_22_207_619;
          st_2 <= `S_2_748;
        end
        `S_2_748: begin
          r2_e0_30_603 <= insn_o_2_1208_0;
          st_2 <= `S_2_749;
        end
        `S_2_749: begin
          r1_e0_25_604 <= r2_e0_30_603;
          st_2 <= `S_2_419;
        end
        `S_2_757: begin
          r3_ror32_2_203_606 <= insn_o_2_1219_0;
          st_2 <= `S_2_760;
        end
        `S_2_760: begin
          r6_ror32_2_204_607 <= insn_o_2_1223_0;
          st_2 <= `S_2_761;
        end
        `S_2_761: begin
          r2_ror32_2_205_608 <= insn_o_2_1225_0;
          st_2 <= `S_2_762;
        end
        `S_2_762: begin
          r1_ror32_2_202_609 <= r2_ror32_2_205_608;
          st_2 <= `S_2_740;
        end
        `S_2_770: begin
          r3_ror32_13_183_611 <= insn_o_2_1236_0;
          st_2 <= `S_2_773;
        end
        `S_2_773: begin
          r6_ror32_13_184_612 <= insn_o_2_1240_0;
          st_2 <= `S_2_774;
        end
        `S_2_774: begin
          r2_ror32_13_185_613 <= insn_o_2_1242_0;
          st_2 <= `S_2_775;
        end
        `S_2_775: begin
          r1_ror32_13_182_614 <= r2_ror32_13_185_613;
          st_2 <= `S_2_743;
        end
        `S_2_783: begin
          r3_ror32_22_208_616 <= insn_o_2_1253_0;
          st_2 <= `S_2_786;
        end
        `S_2_786: begin
          r6_ror32_22_209_617 <= insn_o_2_1257_0;
          st_2 <= `S_2_787;
        end
        `S_2_787: begin
          r2_ror32_22_210_618 <= insn_o_2_1259_0;
          st_2 <= `S_2_788;
        end
        `S_2_788: begin
          r1_ror32_22_207_619 <= r2_ror32_22_210_618;
          st_2 <= `S_2_747;
        end
        `S_2_794: begin
          r5_Maj_11_622 <= insn_o_2_1268_0;
          st_2 <= `S_2_795;
        end
        `S_2_795: begin
          r7_Maj_12_623 <= insn_o_2_1270_0;
          st_2 <= `S_2_796;
        end
        `S_2_796: begin
          r6_Maj_13_625 <= insn_o_2_1272_0;
          st_2 <= `S_2_797;
        end
        `S_2_797: begin
          r4_Maj_14_626 <= insn_o_2_1274_0;
          st_2 <= `S_2_798;
        end
        `S_2_798: begin
          r3_Maj_10_627 <= r4_Maj_14_626;
          st_2 <= `S_2_422;
        end
        `S_2_805: begin
          arg_216_635 <= x_31_628;
          st_2 <= `S_2_823;
        end
        `S_2_806: begin
          r4_e1_33_629 <= r1_ror32_6_217_639;
          st_2 <= `S_2_808;
        end
        `S_2_808: begin
          arg_176_640 <= x_31_628;
          st_2 <= `S_2_836;
        end
        `S_2_809: begin
          r6_e1_34_630 <= r1_ror32_11_177_644;
          st_2 <= `S_2_810;
        end
        `S_2_810: begin
          r3_e1_35_631 <= insn_o_2_1295_0;
          st_2 <= `S_2_812;
        end
        `S_2_812: begin
          arg_211_645 <= x_31_628;
          st_2 <= `S_2_849;
        end
        `S_2_813: begin
          r8_e1_36_632 <= r1_ror32_25_212_649;
          st_2 <= `S_2_814;
        end
        `S_2_814: begin
          r2_e1_37_633 <= insn_o_2_1303_0;
          st_2 <= `S_2_815;
        end
        `S_2_815: begin
          r1_e1_32_634 <= r2_e1_37_633;
          st_2 <= `S_2_431;
        end
        `S_2_823: begin
          r3_ror32_6_218_636 <= insn_o_2_1314_0;
          st_2 <= `S_2_826;
        end
        `S_2_826: begin
          r6_ror32_6_219_637 <= insn_o_2_1318_0;
          st_2 <= `S_2_827;
        end
        `S_2_827: begin
          r2_ror32_6_220_638 <= insn_o_2_1320_0;
          st_2 <= `S_2_828;
        end
        `S_2_828: begin
          r1_ror32_6_217_639 <= r2_ror32_6_220_638;
          st_2 <= `S_2_806;
        end
        `S_2_836: begin
          r3_ror32_11_178_641 <= insn_o_2_1331_0;
          st_2 <= `S_2_839;
        end
        `S_2_839: begin
          r6_ror32_11_179_642 <= insn_o_2_1335_0;
          st_2 <= `S_2_840;
        end
        `S_2_840: begin
          r2_ror32_11_180_643 <= insn_o_2_1337_0;
          st_2 <= `S_2_841;
        end
        `S_2_841: begin
          r1_ror32_11_177_644 <= r2_ror32_11_180_643;
          st_2 <= `S_2_809;
        end
        `S_2_849: begin
          r3_ror32_25_213_646 <= insn_o_2_1348_0;
          st_2 <= `S_2_852;
        end
        `S_2_852: begin
          r6_ror32_25_214_647 <= insn_o_2_1352_0;
          st_2 <= `S_2_853;
        end
        `S_2_853: begin
          r2_ror32_25_215_648 <= insn_o_2_1354_0;
          st_2 <= `S_2_854;
        end
        `S_2_854: begin
          r1_ror32_25_212_649 <= r2_ror32_25_215_648;
          st_2 <= `S_2_813;
        end
        `S_2_860: begin
          r6_Ch_4_652 <= insn_o_2_1363_0;
          st_2 <= `S_2_861;
        end
        `S_2_861: begin
          r5_Ch_5_654 <= insn_o_2_1365_0;
          st_2 <= `S_2_862;
        end
        `S_2_862: begin
          r4_Ch_6_655 <= insn_o_2_1367_0;
          st_2 <= `S_2_863;
        end
        `S_2_863: begin
          r3_Ch_3_656 <= r4_Ch_6_655;
          st_2 <= `S_2_435;
        end
        `S_2_870: begin
          arg_201_664 <= x_24_657;
          st_2 <= `S_2_888;
        end
        `S_2_871: begin
          r4_e0_26_658 <= r1_ror32_2_202_668;
          st_2 <= `S_2_873;
        end
        `S_2_873: begin
          arg_181_669 <= x_24_657;
          st_2 <= `S_2_901;
        end
        `S_2_874: begin
          r6_e0_27_659 <= r1_ror32_13_182_673;
          st_2 <= `S_2_875;
        end
        `S_2_875: begin
          r3_e0_28_660 <= insn_o_2_1388_0;
          st_2 <= `S_2_877;
        end
        `S_2_877: begin
          arg_206_674 <= x_24_657;
          st_2 <= `S_2_914;
        end
        `S_2_878: begin
          r8_e0_29_661 <= r1_ror32_22_207_678;
          st_2 <= `S_2_879;
        end
        `S_2_879: begin
          r2_e0_30_662 <= insn_o_2_1396_0;
          st_2 <= `S_2_880;
        end
        `S_2_880: begin
          r1_e0_25_663 <= r2_e0_30_662;
          st_2 <= `S_2_452;
        end
        `S_2_888: begin
          r3_ror32_2_203_665 <= insn_o_2_1407_0;
          st_2 <= `S_2_891;
        end
        `S_2_891: begin
          r6_ror32_2_204_666 <= insn_o_2_1411_0;
          st_2 <= `S_2_892;
        end
        `S_2_892: begin
          r2_ror32_2_205_667 <= insn_o_2_1413_0;
          st_2 <= `S_2_893;
        end
        `S_2_893: begin
          r1_ror32_2_202_668 <= r2_ror32_2_205_667;
          st_2 <= `S_2_871;
        end
        `S_2_901: begin
          r3_ror32_13_183_670 <= insn_o_2_1424_0;
          st_2 <= `S_2_904;
        end
        `S_2_904: begin
          r6_ror32_13_184_671 <= insn_o_2_1428_0;
          st_2 <= `S_2_905;
        end
        `S_2_905: begin
          r2_ror32_13_185_672 <= insn_o_2_1430_0;
          st_2 <= `S_2_906;
        end
        `S_2_906: begin
          r1_ror32_13_182_673 <= r2_ror32_13_185_672;
          st_2 <= `S_2_874;
        end
        `S_2_914: begin
          r3_ror32_22_208_675 <= insn_o_2_1441_0;
          st_2 <= `S_2_917;
        end
        `S_2_917: begin
          r6_ror32_22_209_676 <= insn_o_2_1445_0;
          st_2 <= `S_2_918;
        end
        `S_2_918: begin
          r2_ror32_22_210_677 <= insn_o_2_1447_0;
          st_2 <= `S_2_919;
        end
        `S_2_919: begin
          r1_ror32_22_207_678 <= r2_ror32_22_210_677;
          st_2 <= `S_2_878;
        end
        `S_2_925: begin
          r5_Maj_11_681 <= insn_o_2_1456_0;
          st_2 <= `S_2_926;
        end
        `S_2_926: begin
          r7_Maj_12_682 <= insn_o_2_1458_0;
          st_2 <= `S_2_927;
        end
        `S_2_927: begin
          r6_Maj_13_684 <= insn_o_2_1460_0;
          st_2 <= `S_2_928;
        end
        `S_2_928: begin
          r4_Maj_14_685 <= insn_o_2_1462_0;
          st_2 <= `S_2_929;
        end
        `S_2_929: begin
          r3_Maj_10_686 <= r4_Maj_14_685;
          st_2 <= `S_2_455;
        end
        `S_2_936: begin
          arg_216_694 <= x_31_687;
          st_2 <= `S_2_954;
        end
        `S_2_937: begin
          r4_e1_33_688 <= r1_ror32_6_217_698;
          st_2 <= `S_2_939;
        end
        `S_2_939: begin
          arg_176_699 <= x_31_687;
          st_2 <= `S_2_967;
        end
        `S_2_940: begin
          r6_e1_34_689 <= r1_ror32_11_177_703;
          st_2 <= `S_2_941;
        end
        `S_2_941: begin
          r3_e1_35_690 <= insn_o_2_1483_0;
          st_2 <= `S_2_943;
        end
        `S_2_943: begin
          arg_211_704 <= x_31_687;
          st_2 <= `S_2_980;
        end
        `S_2_944: begin
          r8_e1_36_691 <= r1_ror32_25_212_708;
          st_2 <= `S_2_945;
        end
        `S_2_945: begin
          r2_e1_37_692 <= insn_o_2_1491_0;
          st_2 <= `S_2_946;
        end
        `S_2_946: begin
          r1_e1_32_693 <= r2_e1_37_692;
          st_2 <= `S_2_464;
        end
        `S_2_954: begin
          r3_ror32_6_218_695 <= insn_o_2_1502_0;
          st_2 <= `S_2_957;
        end
        `S_2_957: begin
          r6_ror32_6_219_696 <= insn_o_2_1506_0;
          st_2 <= `S_2_958;
        end
        `S_2_958: begin
          r2_ror32_6_220_697 <= insn_o_2_1508_0;
          st_2 <= `S_2_959;
        end
        `S_2_959: begin
          r1_ror32_6_217_698 <= r2_ror32_6_220_697;
          st_2 <= `S_2_937;
        end
        `S_2_967: begin
          r3_ror32_11_178_700 <= insn_o_2_1519_0;
          st_2 <= `S_2_970;
        end
        `S_2_970: begin
          r6_ror32_11_179_701 <= insn_o_2_1523_0;
          st_2 <= `S_2_971;
        end
        `S_2_971: begin
          r2_ror32_11_180_702 <= insn_o_2_1525_0;
          st_2 <= `S_2_972;
        end
        `S_2_972: begin
          r1_ror32_11_177_703 <= r2_ror32_11_180_702;
          st_2 <= `S_2_940;
        end
        `S_2_980: begin
          r3_ror32_25_213_705 <= insn_o_2_1536_0;
          st_2 <= `S_2_983;
        end
        `S_2_983: begin
          r6_ror32_25_214_706 <= insn_o_2_1540_0;
          st_2 <= `S_2_984;
        end
        `S_2_984: begin
          r2_ror32_25_215_707 <= insn_o_2_1542_0;
          st_2 <= `S_2_985;
        end
        `S_2_985: begin
          r1_ror32_25_212_708 <= r2_ror32_25_215_707;
          st_2 <= `S_2_944;
        end
        `S_2_991: begin
          r6_Ch_4_711 <= insn_o_2_1551_0;
          st_2 <= `S_2_992;
        end
        `S_2_992: begin
          r5_Ch_5_713 <= insn_o_2_1553_0;
          st_2 <= `S_2_993;
        end
        `S_2_993: begin
          r4_Ch_6_714 <= insn_o_2_1555_0;
          st_2 <= `S_2_994;
        end
        `S_2_994: begin
          r3_Ch_3_715 <= r4_Ch_6_714;
          st_2 <= `S_2_468;
        end
        `S_2_1001: begin
          arg_201_723 <= x_24_716;
          st_2 <= `S_2_1019;
        end
        `S_2_1002: begin
          r4_e0_26_717 <= r1_ror32_2_202_727;
          st_2 <= `S_2_1004;
        end
        `S_2_1004: begin
          arg_181_728 <= x_24_716;
          st_2 <= `S_2_1032;
        end
        `S_2_1005: begin
          r6_e0_27_718 <= r1_ror32_13_182_732;
          st_2 <= `S_2_1006;
        end
        `S_2_1006: begin
          r3_e0_28_719 <= insn_o_2_1576_0;
          st_2 <= `S_2_1008;
        end
        `S_2_1008: begin
          arg_206_733 <= x_24_716;
          st_2 <= `S_2_1045;
        end
        `S_2_1009: begin
          r8_e0_29_720 <= r1_ror32_22_207_737;
          st_2 <= `S_2_1010;
        end
        `S_2_1010: begin
          r2_e0_30_721 <= insn_o_2_1584_0;
          st_2 <= `S_2_1011;
        end
        `S_2_1011: begin
          r1_e0_25_722 <= r2_e0_30_721;
          st_2 <= `S_2_485;
        end
        `S_2_1019: begin
          r3_ror32_2_203_724 <= insn_o_2_1595_0;
          st_2 <= `S_2_1022;
        end
        `S_2_1022: begin
          r6_ror32_2_204_725 <= insn_o_2_1599_0;
          st_2 <= `S_2_1023;
        end
        `S_2_1023: begin
          r2_ror32_2_205_726 <= insn_o_2_1601_0;
          st_2 <= `S_2_1024;
        end
        `S_2_1024: begin
          r1_ror32_2_202_727 <= r2_ror32_2_205_726;
          st_2 <= `S_2_1002;
        end
        `S_2_1032: begin
          r3_ror32_13_183_729 <= insn_o_2_1612_0;
          st_2 <= `S_2_1035;
        end
        `S_2_1035: begin
          r6_ror32_13_184_730 <= insn_o_2_1616_0;
          st_2 <= `S_2_1036;
        end
        `S_2_1036: begin
          r2_ror32_13_185_731 <= insn_o_2_1618_0;
          st_2 <= `S_2_1037;
        end
        `S_2_1037: begin
          r1_ror32_13_182_732 <= r2_ror32_13_185_731;
          st_2 <= `S_2_1005;
        end
        `S_2_1045: begin
          r3_ror32_22_208_734 <= insn_o_2_1629_0;
          st_2 <= `S_2_1048;
        end
        `S_2_1048: begin
          r6_ror32_22_209_735 <= insn_o_2_1633_0;
          st_2 <= `S_2_1049;
        end
        `S_2_1049: begin
          r2_ror32_22_210_736 <= insn_o_2_1635_0;
          st_2 <= `S_2_1050;
        end
        `S_2_1050: begin
          r1_ror32_22_207_737 <= r2_ror32_22_210_736;
          st_2 <= `S_2_1009;
        end
        `S_2_1056: begin
          r5_Maj_11_740 <= insn_o_2_1644_0;
          st_2 <= `S_2_1057;
        end
        `S_2_1057: begin
          r7_Maj_12_741 <= insn_o_2_1646_0;
          st_2 <= `S_2_1058;
        end
        `S_2_1058: begin
          r6_Maj_13_743 <= insn_o_2_1648_0;
          st_2 <= `S_2_1059;
        end
        `S_2_1059: begin
          r4_Maj_14_744 <= insn_o_2_1650_0;
          st_2 <= `S_2_1060;
        end
        `S_2_1060: begin
          r3_Maj_10_745 <= r4_Maj_14_744;
          st_2 <= `S_2_488;
        end
        `S_2_1067: begin
          arg_216_753 <= x_31_746;
          st_2 <= `S_2_1085;
        end
        `S_2_1068: begin
          r4_e1_33_747 <= r1_ror32_6_217_757;
          st_2 <= `S_2_1070;
        end
        `S_2_1070: begin
          arg_176_758 <= x_31_746;
          st_2 <= `S_2_1098;
        end
        `S_2_1071: begin
          r6_e1_34_748 <= r1_ror32_11_177_762;
          st_2 <= `S_2_1072;
        end
        `S_2_1072: begin
          r3_e1_35_749 <= insn_o_2_1671_0;
          st_2 <= `S_2_1074;
        end
        `S_2_1074: begin
          arg_211_763 <= x_31_746;
          st_2 <= `S_2_1111;
        end
        `S_2_1075: begin
          r8_e1_36_750 <= r1_ror32_25_212_767;
          st_2 <= `S_2_1076;
        end
        `S_2_1076: begin
          r2_e1_37_751 <= insn_o_2_1679_0;
          st_2 <= `S_2_1077;
        end
        `S_2_1077: begin
          r1_e1_32_752 <= r2_e1_37_751;
          st_2 <= `S_2_497;
        end
        `S_2_1085: begin
          r3_ror32_6_218_754 <= insn_o_2_1690_0;
          st_2 <= `S_2_1088;
        end
        `S_2_1088: begin
          r6_ror32_6_219_755 <= insn_o_2_1694_0;
          st_2 <= `S_2_1089;
        end
        `S_2_1089: begin
          r2_ror32_6_220_756 <= insn_o_2_1696_0;
          st_2 <= `S_2_1090;
        end
        `S_2_1090: begin
          r1_ror32_6_217_757 <= r2_ror32_6_220_756;
          st_2 <= `S_2_1068;
        end
        `S_2_1098: begin
          r3_ror32_11_178_759 <= insn_o_2_1707_0;
          st_2 <= `S_2_1101;
        end
        `S_2_1101: begin
          r6_ror32_11_179_760 <= insn_o_2_1711_0;
          st_2 <= `S_2_1102;
        end
        `S_2_1102: begin
          r2_ror32_11_180_761 <= insn_o_2_1713_0;
          st_2 <= `S_2_1103;
        end
        `S_2_1103: begin
          r1_ror32_11_177_762 <= r2_ror32_11_180_761;
          st_2 <= `S_2_1071;
        end
        `S_2_1111: begin
          r3_ror32_25_213_764 <= insn_o_2_1724_0;
          st_2 <= `S_2_1114;
        end
        `S_2_1114: begin
          r6_ror32_25_214_765 <= insn_o_2_1728_0;
          st_2 <= `S_2_1115;
        end
        `S_2_1115: begin
          r2_ror32_25_215_766 <= insn_o_2_1730_0;
          st_2 <= `S_2_1116;
        end
        `S_2_1116: begin
          r1_ror32_25_212_767 <= r2_ror32_25_215_766;
          st_2 <= `S_2_1075;
        end
        `S_2_1122: begin
          r6_Ch_4_770 <= insn_o_2_1739_0;
          st_2 <= `S_2_1123;
        end
        `S_2_1123: begin
          r5_Ch_5_772 <= insn_o_2_1741_0;
          st_2 <= `S_2_1124;
        end
        `S_2_1124: begin
          r4_Ch_6_773 <= insn_o_2_1743_0;
          st_2 <= `S_2_1125;
        end
        `S_2_1125: begin
          r3_Ch_3_774 <= r4_Ch_6_773;
          st_2 <= `S_2_501;
        end
        `S_2_1132: begin
          arg_201_782 <= x_24_775;
          st_2 <= `S_2_1150;
        end
        `S_2_1133: begin
          r4_e0_26_776 <= r1_ror32_2_202_786;
          st_2 <= `S_2_1135;
        end
        `S_2_1135: begin
          arg_181_787 <= x_24_775;
          st_2 <= `S_2_1163;
        end
        `S_2_1136: begin
          r6_e0_27_777 <= r1_ror32_13_182_791;
          st_2 <= `S_2_1137;
        end
        `S_2_1137: begin
          r3_e0_28_778 <= insn_o_2_1764_0;
          st_2 <= `S_2_1139;
        end
        `S_2_1139: begin
          arg_206_792 <= x_24_775;
          st_2 <= `S_2_1176;
        end
        `S_2_1140: begin
          r8_e0_29_779 <= r1_ror32_22_207_796;
          st_2 <= `S_2_1141;
        end
        `S_2_1141: begin
          r2_e0_30_780 <= insn_o_2_1772_0;
          st_2 <= `S_2_1142;
        end
        `S_2_1142: begin
          r1_e0_25_781 <= r2_e0_30_780;
          st_2 <= `S_2_518;
        end
        `S_2_1150: begin
          r3_ror32_2_203_783 <= insn_o_2_1783_0;
          st_2 <= `S_2_1153;
        end
        `S_2_1153: begin
          r6_ror32_2_204_784 <= insn_o_2_1787_0;
          st_2 <= `S_2_1154;
        end
        `S_2_1154: begin
          r2_ror32_2_205_785 <= insn_o_2_1789_0;
          st_2 <= `S_2_1155;
        end
        `S_2_1155: begin
          r1_ror32_2_202_786 <= r2_ror32_2_205_785;
          st_2 <= `S_2_1133;
        end
        `S_2_1163: begin
          r3_ror32_13_183_788 <= insn_o_2_1800_0;
          st_2 <= `S_2_1166;
        end
        `S_2_1166: begin
          r6_ror32_13_184_789 <= insn_o_2_1804_0;
          st_2 <= `S_2_1167;
        end
        `S_2_1167: begin
          r2_ror32_13_185_790 <= insn_o_2_1806_0;
          st_2 <= `S_2_1168;
        end
        `S_2_1168: begin
          r1_ror32_13_182_791 <= r2_ror32_13_185_790;
          st_2 <= `S_2_1136;
        end
        `S_2_1176: begin
          r3_ror32_22_208_793 <= insn_o_2_1817_0;
          st_2 <= `S_2_1179;
        end
        `S_2_1179: begin
          r6_ror32_22_209_794 <= insn_o_2_1821_0;
          st_2 <= `S_2_1180;
        end
        `S_2_1180: begin
          r2_ror32_22_210_795 <= insn_o_2_1823_0;
          st_2 <= `S_2_1181;
        end
        `S_2_1181: begin
          r1_ror32_22_207_796 <= r2_ror32_22_210_795;
          st_2 <= `S_2_1140;
        end
        `S_2_1187: begin
          r5_Maj_11_799 <= insn_o_2_1832_0;
          st_2 <= `S_2_1188;
        end
        `S_2_1188: begin
          r7_Maj_12_800 <= insn_o_2_1834_0;
          st_2 <= `S_2_1189;
        end
        `S_2_1189: begin
          r6_Maj_13_802 <= insn_o_2_1836_0;
          st_2 <= `S_2_1190;
        end
        `S_2_1190: begin
          r4_Maj_14_803 <= insn_o_2_1838_0;
          st_2 <= `S_2_1191;
        end
        `S_2_1191: begin
          r3_Maj_10_804 <= r4_Maj_14_803;
          st_2 <= `S_2_521;
        end
        `S_2_1198: begin
          arg_216_812 <= x_31_805;
          st_2 <= `S_2_1216;
        end
        `S_2_1199: begin
          r4_e1_33_806 <= r1_ror32_6_217_816;
          st_2 <= `S_2_1201;
        end
        `S_2_1201: begin
          arg_176_817 <= x_31_805;
          st_2 <= `S_2_1229;
        end
        `S_2_1202: begin
          r6_e1_34_807 <= r1_ror32_11_177_821;
          st_2 <= `S_2_1203;
        end
        `S_2_1203: begin
          r3_e1_35_808 <= insn_o_2_1859_0;
          st_2 <= `S_2_1205;
        end
        `S_2_1205: begin
          arg_211_822 <= x_31_805;
          st_2 <= `S_2_1242;
        end
        `S_2_1206: begin
          r8_e1_36_809 <= r1_ror32_25_212_826;
          st_2 <= `S_2_1207;
        end
        `S_2_1207: begin
          r2_e1_37_810 <= insn_o_2_1867_0;
          st_2 <= `S_2_1208;
        end
        `S_2_1208: begin
          r1_e1_32_811 <= r2_e1_37_810;
          st_2 <= `S_2_530;
        end
        `S_2_1216: begin
          r3_ror32_6_218_813 <= insn_o_2_1878_0;
          st_2 <= `S_2_1219;
        end
        `S_2_1219: begin
          r6_ror32_6_219_814 <= insn_o_2_1882_0;
          st_2 <= `S_2_1220;
        end
        `S_2_1220: begin
          r2_ror32_6_220_815 <= insn_o_2_1884_0;
          st_2 <= `S_2_1221;
        end
        `S_2_1221: begin
          r1_ror32_6_217_816 <= r2_ror32_6_220_815;
          st_2 <= `S_2_1199;
        end
        `S_2_1229: begin
          r3_ror32_11_178_818 <= insn_o_2_1895_0;
          st_2 <= `S_2_1232;
        end
        `S_2_1232: begin
          r6_ror32_11_179_819 <= insn_o_2_1899_0;
          st_2 <= `S_2_1233;
        end
        `S_2_1233: begin
          r2_ror32_11_180_820 <= insn_o_2_1901_0;
          st_2 <= `S_2_1234;
        end
        `S_2_1234: begin
          r1_ror32_11_177_821 <= r2_ror32_11_180_820;
          st_2 <= `S_2_1202;
        end
        `S_2_1242: begin
          r3_ror32_25_213_823 <= insn_o_2_1912_0;
          st_2 <= `S_2_1245;
        end
        `S_2_1245: begin
          r6_ror32_25_214_824 <= insn_o_2_1916_0;
          st_2 <= `S_2_1246;
        end
        `S_2_1246: begin
          r2_ror32_25_215_825 <= insn_o_2_1918_0;
          st_2 <= `S_2_1247;
        end
        `S_2_1247: begin
          r1_ror32_25_212_826 <= r2_ror32_25_215_825;
          st_2 <= `S_2_1206;
        end
        `S_2_1253: begin
          r6_Ch_4_829 <= insn_o_2_1927_0;
          st_2 <= `S_2_1254;
        end
        `S_2_1254: begin
          r5_Ch_5_831 <= insn_o_2_1929_0;
          st_2 <= `S_2_1255;
        end
        `S_2_1255: begin
          r4_Ch_6_832 <= insn_o_2_1931_0;
          st_2 <= `S_2_1256;
        end
        `S_2_1256: begin
          r3_Ch_3_833 <= r4_Ch_6_832;
          st_2 <= `S_2_534;
        end
        `S_2_1263: begin
          arg_201_841 <= x_24_834;
          st_2 <= `S_2_1281;
        end
        `S_2_1264: begin
          r4_e0_26_835 <= r1_ror32_2_202_845;
          st_2 <= `S_2_1266;
        end
        `S_2_1266: begin
          arg_181_846 <= x_24_834;
          st_2 <= `S_2_1294;
        end
        `S_2_1267: begin
          r6_e0_27_836 <= r1_ror32_13_182_850;
          st_2 <= `S_2_1268;
        end
        `S_2_1268: begin
          r3_e0_28_837 <= insn_o_2_1952_0;
          st_2 <= `S_2_1270;
        end
        `S_2_1270: begin
          arg_206_851 <= x_24_834;
          st_2 <= `S_2_1307;
        end
        `S_2_1271: begin
          r8_e0_29_838 <= r1_ror32_22_207_855;
          st_2 <= `S_2_1272;
        end
        `S_2_1272: begin
          r2_e0_30_839 <= insn_o_2_1960_0;
          st_2 <= `S_2_1273;
        end
        `S_2_1273: begin
          r1_e0_25_840 <= r2_e0_30_839;
          st_2 <= `S_2_551;
        end
        `S_2_1281: begin
          r3_ror32_2_203_842 <= insn_o_2_1971_0;
          st_2 <= `S_2_1284;
        end
        `S_2_1284: begin
          r6_ror32_2_204_843 <= insn_o_2_1975_0;
          st_2 <= `S_2_1285;
        end
        `S_2_1285: begin
          r2_ror32_2_205_844 <= insn_o_2_1977_0;
          st_2 <= `S_2_1286;
        end
        `S_2_1286: begin
          r1_ror32_2_202_845 <= r2_ror32_2_205_844;
          st_2 <= `S_2_1264;
        end
        `S_2_1294: begin
          r3_ror32_13_183_847 <= insn_o_2_1988_0;
          st_2 <= `S_2_1297;
        end
        `S_2_1297: begin
          r6_ror32_13_184_848 <= insn_o_2_1992_0;
          st_2 <= `S_2_1298;
        end
        `S_2_1298: begin
          r2_ror32_13_185_849 <= insn_o_2_1994_0;
          st_2 <= `S_2_1299;
        end
        `S_2_1299: begin
          r1_ror32_13_182_850 <= r2_ror32_13_185_849;
          st_2 <= `S_2_1267;
        end
        `S_2_1307: begin
          r3_ror32_22_208_852 <= insn_o_2_2005_0;
          st_2 <= `S_2_1310;
        end
        `S_2_1310: begin
          r6_ror32_22_209_853 <= insn_o_2_2009_0;
          st_2 <= `S_2_1311;
        end
        `S_2_1311: begin
          r2_ror32_22_210_854 <= insn_o_2_2011_0;
          st_2 <= `S_2_1312;
        end
        `S_2_1312: begin
          r1_ror32_22_207_855 <= r2_ror32_22_210_854;
          st_2 <= `S_2_1271;
        end
        `S_2_1318: begin
          r5_Maj_11_858 <= insn_o_2_2020_0;
          st_2 <= `S_2_1319;
        end
        `S_2_1319: begin
          r7_Maj_12_859 <= insn_o_2_2022_0;
          st_2 <= `S_2_1320;
        end
        `S_2_1320: begin
          r6_Maj_13_861 <= insn_o_2_2024_0;
          st_2 <= `S_2_1321;
        end
        `S_2_1321: begin
          r4_Maj_14_862 <= insn_o_2_2026_0;
          st_2 <= `S_2_1322;
        end
        `S_2_1322: begin
          r3_Maj_10_863 <= r4_Maj_14_862;
          st_2 <= `S_2_554;
        end
        `S_2_1329: begin
          arg_216_871 <= x_31_864;
          st_2 <= `S_2_1347;
        end
        `S_2_1330: begin
          r4_e1_33_865 <= r1_ror32_6_217_875;
          st_2 <= `S_2_1332;
        end
        `S_2_1332: begin
          arg_176_876 <= x_31_864;
          st_2 <= `S_2_1360;
        end
        `S_2_1333: begin
          r6_e1_34_866 <= r1_ror32_11_177_880;
          st_2 <= `S_2_1334;
        end
        `S_2_1334: begin
          r3_e1_35_867 <= insn_o_2_2047_0;
          st_2 <= `S_2_1336;
        end
        `S_2_1336: begin
          arg_211_881 <= x_31_864;
          st_2 <= `S_2_1373;
        end
        `S_2_1337: begin
          r8_e1_36_868 <= r1_ror32_25_212_885;
          st_2 <= `S_2_1338;
        end
        `S_2_1338: begin
          r2_e1_37_869 <= insn_o_2_2055_0;
          st_2 <= `S_2_1339;
        end
        `S_2_1339: begin
          r1_e1_32_870 <= r2_e1_37_869;
          st_2 <= `S_2_563;
        end
        `S_2_1347: begin
          r3_ror32_6_218_872 <= insn_o_2_2066_0;
          st_2 <= `S_2_1350;
        end
        `S_2_1350: begin
          r6_ror32_6_219_873 <= insn_o_2_2070_0;
          st_2 <= `S_2_1351;
        end
        `S_2_1351: begin
          r2_ror32_6_220_874 <= insn_o_2_2072_0;
          st_2 <= `S_2_1352;
        end
        `S_2_1352: begin
          r1_ror32_6_217_875 <= r2_ror32_6_220_874;
          st_2 <= `S_2_1330;
        end
        `S_2_1360: begin
          r3_ror32_11_178_877 <= insn_o_2_2083_0;
          st_2 <= `S_2_1363;
        end
        `S_2_1363: begin
          r6_ror32_11_179_878 <= insn_o_2_2087_0;
          st_2 <= `S_2_1364;
        end
        `S_2_1364: begin
          r2_ror32_11_180_879 <= insn_o_2_2089_0;
          st_2 <= `S_2_1365;
        end
        `S_2_1365: begin
          r1_ror32_11_177_880 <= r2_ror32_11_180_879;
          st_2 <= `S_2_1333;
        end
        `S_2_1373: begin
          r3_ror32_25_213_882 <= insn_o_2_2100_0;
          st_2 <= `S_2_1376;
        end
        `S_2_1376: begin
          r6_ror32_25_214_883 <= insn_o_2_2104_0;
          st_2 <= `S_2_1377;
        end
        `S_2_1377: begin
          r2_ror32_25_215_884 <= insn_o_2_2106_0;
          st_2 <= `S_2_1378;
        end
        `S_2_1378: begin
          r1_ror32_25_212_885 <= r2_ror32_25_215_884;
          st_2 <= `S_2_1337;
        end
        `S_2_1384: begin
          r6_Ch_4_888 <= insn_o_2_2115_0;
          st_2 <= `S_2_1385;
        end
        `S_2_1385: begin
          r5_Ch_5_890 <= insn_o_2_2117_0;
          st_2 <= `S_2_1386;
        end
        `S_2_1386: begin
          r4_Ch_6_891 <= insn_o_2_2119_0;
          st_2 <= `S_2_1387;
        end
        `S_2_1387: begin
          r3_Ch_3_892 <= r4_Ch_6_891;
          st_2 <= `S_2_567;
        end
        `S_2_1394: begin
          arg_201_900 <= x_24_893;
          st_2 <= `S_2_1412;
        end
        `S_2_1395: begin
          r4_e0_26_894 <= r1_ror32_2_202_904;
          st_2 <= `S_2_1397;
        end
        `S_2_1397: begin
          arg_181_905 <= x_24_893;
          st_2 <= `S_2_1425;
        end
        `S_2_1398: begin
          r6_e0_27_895 <= r1_ror32_13_182_909;
          st_2 <= `S_2_1399;
        end
        `S_2_1399: begin
          r3_e0_28_896 <= insn_o_2_2140_0;
          st_2 <= `S_2_1401;
        end
        `S_2_1401: begin
          arg_206_910 <= x_24_893;
          st_2 <= `S_2_1438;
        end
        `S_2_1402: begin
          r8_e0_29_897 <= r1_ror32_22_207_914;
          st_2 <= `S_2_1403;
        end
        `S_2_1403: begin
          r2_e0_30_898 <= insn_o_2_2148_0;
          st_2 <= `S_2_1404;
        end
        `S_2_1404: begin
          r1_e0_25_899 <= r2_e0_30_898;
          st_2 <= `S_2_584;
        end
        `S_2_1412: begin
          r3_ror32_2_203_901 <= insn_o_2_2159_0;
          st_2 <= `S_2_1415;
        end
        `S_2_1415: begin
          r6_ror32_2_204_902 <= insn_o_2_2163_0;
          st_2 <= `S_2_1416;
        end
        `S_2_1416: begin
          r2_ror32_2_205_903 <= insn_o_2_2165_0;
          st_2 <= `S_2_1417;
        end
        `S_2_1417: begin
          r1_ror32_2_202_904 <= r2_ror32_2_205_903;
          st_2 <= `S_2_1395;
        end
        `S_2_1425: begin
          r3_ror32_13_183_906 <= insn_o_2_2176_0;
          st_2 <= `S_2_1428;
        end
        `S_2_1428: begin
          r6_ror32_13_184_907 <= insn_o_2_2180_0;
          st_2 <= `S_2_1429;
        end
        `S_2_1429: begin
          r2_ror32_13_185_908 <= insn_o_2_2182_0;
          st_2 <= `S_2_1430;
        end
        `S_2_1430: begin
          r1_ror32_13_182_909 <= r2_ror32_13_185_908;
          st_2 <= `S_2_1398;
        end
        `S_2_1438: begin
          r3_ror32_22_208_911 <= insn_o_2_2193_0;
          st_2 <= `S_2_1441;
        end
        `S_2_1441: begin
          r6_ror32_22_209_912 <= insn_o_2_2197_0;
          st_2 <= `S_2_1442;
        end
        `S_2_1442: begin
          r2_ror32_22_210_913 <= insn_o_2_2199_0;
          st_2 <= `S_2_1443;
        end
        `S_2_1443: begin
          r1_ror32_22_207_914 <= r2_ror32_22_210_913;
          st_2 <= `S_2_1402;
        end
        `S_2_1449: begin
          r5_Maj_11_917 <= insn_o_2_2208_0;
          st_2 <= `S_2_1450;
        end
        `S_2_1450: begin
          r7_Maj_12_918 <= insn_o_2_2210_0;
          st_2 <= `S_2_1451;
        end
        `S_2_1451: begin
          r6_Maj_13_920 <= insn_o_2_2212_0;
          st_2 <= `S_2_1452;
        end
        `S_2_1452: begin
          r4_Maj_14_921 <= insn_o_2_2214_0;
          st_2 <= `S_2_1453;
        end
        `S_2_1453: begin
          r3_Maj_10_922 <= r4_Maj_14_921;
          st_2 <= `S_2_587;
        end
        `S_2_1460: begin
          arg_216_930 <= x_31_923;
          st_2 <= `S_2_1478;
        end
        `S_2_1461: begin
          r4_e1_33_924 <= r1_ror32_6_217_934;
          st_2 <= `S_2_1463;
        end
        `S_2_1463: begin
          arg_176_935 <= x_31_923;
          st_2 <= `S_2_1491;
        end
        `S_2_1464: begin
          r6_e1_34_925 <= r1_ror32_11_177_939;
          st_2 <= `S_2_1465;
        end
        `S_2_1465: begin
          r3_e1_35_926 <= insn_o_2_2235_0;
          st_2 <= `S_2_1467;
        end
        `S_2_1467: begin
          arg_211_940 <= x_31_923;
          st_2 <= `S_2_1504;
        end
        `S_2_1468: begin
          r8_e1_36_927 <= r1_ror32_25_212_944;
          st_2 <= `S_2_1469;
        end
        `S_2_1469: begin
          r2_e1_37_928 <= insn_o_2_2243_0;
          st_2 <= `S_2_1470;
        end
        `S_2_1470: begin
          r1_e1_32_929 <= r2_e1_37_928;
          st_2 <= `S_2_596;
        end
        `S_2_1478: begin
          r3_ror32_6_218_931 <= insn_o_2_2254_0;
          st_2 <= `S_2_1481;
        end
        `S_2_1481: begin
          r6_ror32_6_219_932 <= insn_o_2_2258_0;
          st_2 <= `S_2_1482;
        end
        `S_2_1482: begin
          r2_ror32_6_220_933 <= insn_o_2_2260_0;
          st_2 <= `S_2_1483;
        end
        `S_2_1483: begin
          r1_ror32_6_217_934 <= r2_ror32_6_220_933;
          st_2 <= `S_2_1461;
        end
        `S_2_1491: begin
          r3_ror32_11_178_936 <= insn_o_2_2271_0;
          st_2 <= `S_2_1494;
        end
        `S_2_1494: begin
          r6_ror32_11_179_937 <= insn_o_2_2275_0;
          st_2 <= `S_2_1495;
        end
        `S_2_1495: begin
          r2_ror32_11_180_938 <= insn_o_2_2277_0;
          st_2 <= `S_2_1496;
        end
        `S_2_1496: begin
          r1_ror32_11_177_939 <= r2_ror32_11_180_938;
          st_2 <= `S_2_1464;
        end
        `S_2_1504: begin
          r3_ror32_25_213_941 <= insn_o_2_2288_0;
          st_2 <= `S_2_1507;
        end
        `S_2_1507: begin
          r6_ror32_25_214_942 <= insn_o_2_2292_0;
          st_2 <= `S_2_1508;
        end
        `S_2_1508: begin
          r2_ror32_25_215_943 <= insn_o_2_2294_0;
          st_2 <= `S_2_1509;
        end
        `S_2_1509: begin
          r1_ror32_25_212_944 <= r2_ror32_25_215_943;
          st_2 <= `S_2_1468;
        end
        `S_2_1515: begin
          r6_Ch_4_947 <= insn_o_2_2303_0;
          st_2 <= `S_2_1516;
        end
        `S_2_1516: begin
          r5_Ch_5_949 <= insn_o_2_2305_0;
          st_2 <= `S_2_1517;
        end
        `S_2_1517: begin
          r4_Ch_6_950 <= insn_o_2_2307_0;
          st_2 <= `S_2_1518;
        end
        `S_2_1518: begin
          r3_Ch_3_951 <= r4_Ch_6_950;
          st_2 <= `S_2_600;
        end
        `S_2_1525: begin
          arg_201_959 <= x_24_952;
          st_2 <= `S_2_1543;
        end
        `S_2_1526: begin
          r4_e0_26_953 <= r1_ror32_2_202_963;
          st_2 <= `S_2_1528;
        end
        `S_2_1528: begin
          arg_181_964 <= x_24_952;
          st_2 <= `S_2_1556;
        end
        `S_2_1529: begin
          r6_e0_27_954 <= r1_ror32_13_182_968;
          st_2 <= `S_2_1530;
        end
        `S_2_1530: begin
          r3_e0_28_955 <= insn_o_2_2328_0;
          st_2 <= `S_2_1532;
        end
        `S_2_1532: begin
          arg_206_969 <= x_24_952;
          st_2 <= `S_2_1569;
        end
        `S_2_1533: begin
          r8_e0_29_956 <= r1_ror32_22_207_973;
          st_2 <= `S_2_1534;
        end
        `S_2_1534: begin
          r2_e0_30_957 <= insn_o_2_2336_0;
          st_2 <= `S_2_1535;
        end
        `S_2_1535: begin
          r1_e0_25_958 <= r2_e0_30_957;
          st_2 <= `S_2_617;
        end
        `S_2_1543: begin
          r3_ror32_2_203_960 <= insn_o_2_2347_0;
          st_2 <= `S_2_1546;
        end
        `S_2_1546: begin
          r6_ror32_2_204_961 <= insn_o_2_2351_0;
          st_2 <= `S_2_1547;
        end
        `S_2_1547: begin
          r2_ror32_2_205_962 <= insn_o_2_2353_0;
          st_2 <= `S_2_1548;
        end
        `S_2_1548: begin
          r1_ror32_2_202_963 <= r2_ror32_2_205_962;
          st_2 <= `S_2_1526;
        end
        `S_2_1556: begin
          r3_ror32_13_183_965 <= insn_o_2_2364_0;
          st_2 <= `S_2_1559;
        end
        `S_2_1559: begin
          r6_ror32_13_184_966 <= insn_o_2_2368_0;
          st_2 <= `S_2_1560;
        end
        `S_2_1560: begin
          r2_ror32_13_185_967 <= insn_o_2_2370_0;
          st_2 <= `S_2_1561;
        end
        `S_2_1561: begin
          r1_ror32_13_182_968 <= r2_ror32_13_185_967;
          st_2 <= `S_2_1529;
        end
        `S_2_1569: begin
          r3_ror32_22_208_970 <= insn_o_2_2381_0;
          st_2 <= `S_2_1572;
        end
        `S_2_1572: begin
          r6_ror32_22_209_971 <= insn_o_2_2385_0;
          st_2 <= `S_2_1573;
        end
        `S_2_1573: begin
          r2_ror32_22_210_972 <= insn_o_2_2387_0;
          st_2 <= `S_2_1574;
        end
        `S_2_1574: begin
          r1_ror32_22_207_973 <= r2_ror32_22_210_972;
          st_2 <= `S_2_1533;
        end
        `S_2_1580: begin
          r5_Maj_11_976 <= insn_o_2_2396_0;
          st_2 <= `S_2_1581;
        end
        `S_2_1581: begin
          r7_Maj_12_977 <= insn_o_2_2398_0;
          st_2 <= `S_2_1582;
        end
        `S_2_1582: begin
          r6_Maj_13_979 <= insn_o_2_2400_0;
          st_2 <= `S_2_1583;
        end
        `S_2_1583: begin
          r4_Maj_14_980 <= insn_o_2_2402_0;
          st_2 <= `S_2_1584;
        end
        `S_2_1584: begin
          r3_Maj_10_981 <= r4_Maj_14_980;
          st_2 <= `S_2_620;
        end
        `S_2_1591: begin
          arg_216_989 <= x_31_982;
          st_2 <= `S_2_1609;
        end
        `S_2_1592: begin
          r4_e1_33_983 <= r1_ror32_6_217_993;
          st_2 <= `S_2_1594;
        end
        `S_2_1594: begin
          arg_176_994 <= x_31_982;
          st_2 <= `S_2_1622;
        end
        `S_2_1595: begin
          r6_e1_34_984 <= r1_ror32_11_177_998;
          st_2 <= `S_2_1596;
        end
        `S_2_1596: begin
          r3_e1_35_985 <= insn_o_2_2423_0;
          st_2 <= `S_2_1598;
        end
        `S_2_1598: begin
          arg_211_999 <= x_31_982;
          st_2 <= `S_2_1635;
        end
        `S_2_1599: begin
          r8_e1_36_986 <= r1_ror32_25_212_1003;
          st_2 <= `S_2_1600;
        end
        `S_2_1600: begin
          r2_e1_37_987 <= insn_o_2_2431_0;
          st_2 <= `S_2_1601;
        end
        `S_2_1601: begin
          r1_e1_32_988 <= r2_e1_37_987;
          st_2 <= `S_2_629;
        end
        `S_2_1609: begin
          r3_ror32_6_218_990 <= insn_o_2_2442_0;
          st_2 <= `S_2_1612;
        end
        `S_2_1612: begin
          r6_ror32_6_219_991 <= insn_o_2_2446_0;
          st_2 <= `S_2_1613;
        end
        `S_2_1613: begin
          r2_ror32_6_220_992 <= insn_o_2_2448_0;
          st_2 <= `S_2_1614;
        end
        `S_2_1614: begin
          r1_ror32_6_217_993 <= r2_ror32_6_220_992;
          st_2 <= `S_2_1592;
        end
        `S_2_1622: begin
          r3_ror32_11_178_995 <= insn_o_2_2459_0;
          st_2 <= `S_2_1625;
        end
        `S_2_1625: begin
          r6_ror32_11_179_996 <= insn_o_2_2463_0;
          st_2 <= `S_2_1626;
        end
        `S_2_1626: begin
          r2_ror32_11_180_997 <= insn_o_2_2465_0;
          st_2 <= `S_2_1627;
        end
        `S_2_1627: begin
          r1_ror32_11_177_998 <= r2_ror32_11_180_997;
          st_2 <= `S_2_1595;
        end
        `S_2_1635: begin
          r3_ror32_25_213_1000 <= insn_o_2_2476_0;
          st_2 <= `S_2_1638;
        end
        `S_2_1638: begin
          r6_ror32_25_214_1001 <= insn_o_2_2480_0;
          st_2 <= `S_2_1639;
        end
        `S_2_1639: begin
          r2_ror32_25_215_1002 <= insn_o_2_2482_0;
          st_2 <= `S_2_1640;
        end
        `S_2_1640: begin
          r1_ror32_25_212_1003 <= r2_ror32_25_215_1002;
          st_2 <= `S_2_1599;
        end
        `S_2_1646: begin
          r6_Ch_4_1006 <= insn_o_2_2491_0;
          st_2 <= `S_2_1647;
        end
        `S_2_1647: begin
          r5_Ch_5_1008 <= insn_o_2_2493_0;
          st_2 <= `S_2_1648;
        end
        `S_2_1648: begin
          r4_Ch_6_1009 <= insn_o_2_2495_0;
          st_2 <= `S_2_1649;
        end
        `S_2_1649: begin
          r3_Ch_3_1010 <= r4_Ch_6_1009;
          st_2 <= `S_2_633;
        end
        `S_2_1656: begin
          arg_201_1018 <= x_24_1011;
          st_2 <= `S_2_1674;
        end
        `S_2_1657: begin
          r4_e0_26_1012 <= r1_ror32_2_202_1022;
          st_2 <= `S_2_1659;
        end
        `S_2_1659: begin
          arg_181_1023 <= x_24_1011;
          st_2 <= `S_2_1687;
        end
        `S_2_1660: begin
          r6_e0_27_1013 <= r1_ror32_13_182_1027;
          st_2 <= `S_2_1661;
        end
        `S_2_1661: begin
          r3_e0_28_1014 <= insn_o_2_2516_0;
          st_2 <= `S_2_1663;
        end
        `S_2_1663: begin
          arg_206_1028 <= x_24_1011;
          st_2 <= `S_2_1700;
        end
        `S_2_1664: begin
          r8_e0_29_1015 <= r1_ror32_22_207_1032;
          st_2 <= `S_2_1665;
        end
        `S_2_1665: begin
          r2_e0_30_1016 <= insn_o_2_2524_0;
          st_2 <= `S_2_1666;
        end
        `S_2_1666: begin
          r1_e0_25_1017 <= r2_e0_30_1016;
          st_2 <= `S_2_650;
        end
        `S_2_1674: begin
          r3_ror32_2_203_1019 <= insn_o_2_2535_0;
          st_2 <= `S_2_1677;
        end
        `S_2_1677: begin
          r6_ror32_2_204_1020 <= insn_o_2_2539_0;
          st_2 <= `S_2_1678;
        end
        `S_2_1678: begin
          r2_ror32_2_205_1021 <= insn_o_2_2541_0;
          st_2 <= `S_2_1679;
        end
        `S_2_1679: begin
          r1_ror32_2_202_1022 <= r2_ror32_2_205_1021;
          st_2 <= `S_2_1657;
        end
        `S_2_1687: begin
          r3_ror32_13_183_1024 <= insn_o_2_2552_0;
          st_2 <= `S_2_1690;
        end
        `S_2_1690: begin
          r6_ror32_13_184_1025 <= insn_o_2_2556_0;
          st_2 <= `S_2_1691;
        end
        `S_2_1691: begin
          r2_ror32_13_185_1026 <= insn_o_2_2558_0;
          st_2 <= `S_2_1692;
        end
        `S_2_1692: begin
          r1_ror32_13_182_1027 <= r2_ror32_13_185_1026;
          st_2 <= `S_2_1660;
        end
        `S_2_1700: begin
          r3_ror32_22_208_1029 <= insn_o_2_2569_0;
          st_2 <= `S_2_1703;
        end
        `S_2_1703: begin
          r6_ror32_22_209_1030 <= insn_o_2_2573_0;
          st_2 <= `S_2_1704;
        end
        `S_2_1704: begin
          r2_ror32_22_210_1031 <= insn_o_2_2575_0;
          st_2 <= `S_2_1705;
        end
        `S_2_1705: begin
          r1_ror32_22_207_1032 <= r2_ror32_22_210_1031;
          st_2 <= `S_2_1664;
        end
        `S_2_1711: begin
          r5_Maj_11_1035 <= insn_o_2_2584_0;
          st_2 <= `S_2_1712;
        end
        `S_2_1712: begin
          r7_Maj_12_1036 <= insn_o_2_2586_0;
          st_2 <= `S_2_1713;
        end
        `S_2_1713: begin
          r6_Maj_13_1038 <= insn_o_2_2588_0;
          st_2 <= `S_2_1714;
        end
        `S_2_1714: begin
          r4_Maj_14_1039 <= insn_o_2_2590_0;
          st_2 <= `S_2_1715;
        end
        `S_2_1715: begin
          r3_Maj_10_1040 <= r4_Maj_14_1039;
          st_2 <= `S_2_653;
        end
      endcase
    end
  end
  SRAM_4_32_2 SRAM_4_32_2_inst_2_15(.clk(clk), .rst(rst), .addr_0_i(mem_1_2_15_p0_addr), .rdata_0_o(mem_1_2_15_p0_rdata), .wdata_0_i(mem_1_2_15_p0_wdata), .write_en_0_i(mem_1_2_15_p0_wen), .addr_1_i(mem_1_2_15_p1_addr), .rdata_1_o(mem_1_2_15_p1_rdata), .wdata_1_i(mem_1_2_15_p1_wdata), .write_en_1_i(mem_1_2_15_p1_wen));
  axi_master_controller_a4rd32 inst_2_16_axi_master_controller_a4rd32(.clk(clk), .rst(rst), .sram_addr(mem_1_2_15_p1_addr), .sram_wdata(mem_1_2_15_p1_wdata), .sram_rdata(mem_1_2_15_p1_rdata), .sram_wen(mem_1_2_15_p1_wen), .sram_EXCLUSIVE(1), .sram_req(/*not connected*/), .sram_ack(1), .addr(axi_addr2_16), .wen(axi_wen2_16), .req(axi_req2_16), .len(axi_len2_16), .start(axi_start2_16), .ack(axi_ack2_16) , .ARADDR(buf_ARADDR), .ARVALID(buf_ARVALID), .ARREADY(buf_ARREADY), .ARLEN(buf_ARLEN), .ARSIZE(buf_ARSIZE), .RVALID(buf_RVALID), .RDATA(buf_RDATA), .RREADY(buf_RREADY), .RLAST(buf_RLAST), .AWADDR(buf_AWADDR), .AWVALID(buf_AWVALID), .AWREADY(buf_AWREADY), .AWLEN(buf_AWLEN), .AWSIZE(buf_AWSIZE), .WVALID(buf_WVALID), .WREADY(buf_WREADY), .WDATA(buf_WDATA), .WLAST(buf_WLAST), .BVALID(buf_BVALID), .BREADY(buf_BREADY), .BRESP(buf_BRESP));
  SRAM_3_32 SRAM_3_32_inst_2(.clk(clk), .rst(rst), .addr_i(sram_addr_2), .rdata_o(sram_rdata_2), .wdata_i(sram_wdata_2), .write_en_i(sram_wdata_en_2));
  SRAM_6_32 SRAM_6_32_inst_20(.clk(clk), .rst(rst), .addr_i(sram_addr_20), .rdata_o(sram_rdata_20), .wdata_i(sram_wdata_20), .write_en_i(sram_wdata_en_20));
  SRAM_6_32 SRAM_6_32_inst_21(.clk(clk), .rst(rst), .addr_i(sram_addr_21), .rdata_o(sram_rdata_21), .wdata_i(sram_wdata_21), .write_en_i(sram_wdata_en_21));

endmodule // main
module sha256(clk, rst, buf_ARADDR, buf_ARVALID, buf_ARREADY, buf_ARLEN, buf_ARSIZE, buf_RVALID, buf_RDATA, buf_RREADY, buf_RLAST, buf_AWADDR, buf_AWVALID, buf_AWREADY, buf_AWLEN, buf_AWSIZE, buf_WVALID, buf_WREADY, buf_WDATA, buf_WLAST, buf_BVALID, buf_BREADY, buf_BRESP, sha256_req_valid, sha256_req_ready, sha256_req_busy, sha256_res_valid, sha256_res_ready, sha256_req_0, sha256_req_1, sha256_res_0);
  input clk;
  input rst;
  output [31:0] buf_ARADDR;
  output buf_ARVALID;
  input buf_ARREADY;
  output [7:0] buf_ARLEN;
  output [2:0] buf_ARSIZE;
  input buf_RVALID;
  input [31:0] buf_RDATA;
  output buf_RREADY;
  input buf_RLAST;
  output [31:0] buf_AWADDR;
  output buf_AWVALID;
  input buf_AWREADY;
  output [7:0] buf_AWLEN;
  output [2:0] buf_AWSIZE;
  output buf_WVALID;
  input buf_WREADY;
  output [31:0] buf_WDATA;
  output buf_WLAST;
  input buf_BVALID;
  output buf_BREADY;
  input [1:0] buf_BRESP;
  input sha256_req_valid;
  output sha256_req_ready;
  output sha256_req_busy;
  output sha256_res_valid;
  input sha256_res_ready;
  input [31:0] sha256_req_0;
  input [31:0] sha256_req_1;
  output [255:0] sha256_res_0;
  main main_inst(.clk(clk), .rst(rst), .buf_ARADDR(buf_ARADDR), .buf_ARVALID(buf_ARVALID), .buf_ARREADY(buf_ARREADY), .buf_ARLEN(buf_ARLEN), .buf_ARSIZE(buf_ARSIZE), .buf_RVALID(buf_RVALID), .buf_RDATA(buf_RDATA), .buf_RREADY(buf_RREADY), .buf_RLAST(buf_RLAST), .buf_AWADDR(buf_AWADDR), .buf_AWVALID(buf_AWVALID), .buf_AWREADY(buf_AWREADY), .buf_AWLEN(buf_AWLEN), .buf_AWSIZE(buf_AWSIZE), .buf_WVALID(buf_WVALID), .buf_WREADY(buf_WREADY), .buf_WDATA(buf_WDATA), .buf_WLAST(buf_WLAST), .buf_BVALID(buf_BVALID), .buf_BREADY(buf_BREADY), .buf_BRESP(buf_BRESP), .sha256_req_valid(sha256_req_valid), .sha256_req_ready(sha256_req_ready), .sha256_req_busy(sha256_req_busy), .sha256_res_valid(sha256_res_valid), .sha256_res_ready(sha256_res_ready), .sha256_req_0(sha256_req_0), .sha256_req_1(sha256_req_1), .sha256_res_0(sha256_res_0));
endmodule
