// Generated from iroha-0.0.1.

// SRAM(2 port(s))
module SRAM_4_32_2(clk, rst, addr_0_i, rdata_0_o, wdata_0_i, write_en_0_i, addr_1_i, rdata_1_o, wdata_1_i, write_en_1_i);
  input clk;
  input rst;
  input [3:0] addr_0_i;
  output [31:0] rdata_0_o;
  input [31:0] wdata_0_i;
  input write_en_0_i;

  reg [31:0] rdata_0_o;

  input [3:0] addr_1_i;
  output [31:0] rdata_1_o;
  input [31:0] wdata_1_i;
  input write_en_1_i;

  reg [31:0] rdata_1_o;

  reg [31:0] data [0:15];

  always @(posedge clk) begin
    if (rst) begin
    end else begin
      if (write_en_0_i) begin
        data[addr_0_i] <= wdata_0_i;
      end
      if (write_en_1_i) begin
        data[addr_1_i] <= wdata_1_i;
      end
    end
  end
  // Read
  always @(addr_0_i or clk) begin
    rdata_0_o = data[addr_0_i];
  end
  always @(addr_1_i or clk) begin
    rdata_1_o = data[addr_1_i];
  end
endmodule


// SRAM(1 port(s))
module SRAM_3_32(clk, rst, addr_i, rdata_o, wdata_i, write_en_i);
  input clk;
  input rst;
  input [2:0] addr_i;
  output [31:0] rdata_o;
  input [31:0] wdata_i;
  input write_en_i;

  reg [31:0] rdata_o;

  reg [31:0] data [0:7];

  always @(posedge clk) begin
    if (rst) begin
      data[0] <= 0;
      data[1] <= 0;
      data[2] <= 0;
      data[3] <= 0;
      data[4] <= 0;
      data[5] <= 0;
      data[6] <= 0;
      data[7] <= 0;
    end else begin
      if (write_en_i) begin
        data[addr_i] <= wdata_i;
      end
    end
  end
  // Read
  always @(addr_i or clk) begin
    rdata_o = data[addr_i];
  end
endmodule


// SRAM(1 port(s))
module SRAM_6_32(clk, rst, addr_i, rdata_o, wdata_i, write_en_i);
  input clk;
  input rst;
  input [5:0] addr_i;
  output [31:0] rdata_o;
  input [31:0] wdata_i;
  input write_en_i;

  reg [31:0] rdata_o;

  reg [31:0] data [0:63];

  always @(posedge clk) begin
    if (rst) begin
      data[0] <= 1116352408;
      data[1] <= 1899447441;
      data[2] <= -1245643825;
      data[3] <= -373957723;
      data[4] <= 961987163;
      data[5] <= 1508970993;
      data[6] <= -1841331548;
      data[7] <= -1424204075;
      data[8] <= -670586216;
      data[9] <= 310598401;
      data[10] <= 607225278;
      data[11] <= 1426881987;
      data[12] <= 1925078388;
      data[13] <= -2132889090;
      data[14] <= -1680079193;
      data[15] <= -1046744716;
      data[16] <= -459576895;
      data[17] <= -272742522;
      data[18] <= 264347078;
      data[19] <= 604807628;
      data[20] <= 770255983;
      data[21] <= 1249150122;
      data[22] <= 1555081692;
      data[23] <= 1996064986;
      data[24] <= -1740746414;
      data[25] <= -1473132947;
      data[26] <= -1341970488;
      data[27] <= -1084653625;
      data[28] <= -958395405;
      data[29] <= -710438585;
      data[30] <= 113926993;
      data[31] <= 338241895;
      data[32] <= 666307205;
      data[33] <= 773529912;
      data[34] <= 1294757372;
      data[35] <= 1396182291;
      data[36] <= 1695183700;
      data[37] <= 1986661051;
      data[38] <= -2117940946;
      data[39] <= -1838011259;
      data[40] <= -1564481375;
      data[41] <= -1474664885;
      data[42] <= -1035236496;
      data[43] <= -949202525;
      data[44] <= -778901479;
      data[45] <= -694614492;
      data[46] <= -200395387;
      data[47] <= 275423344;
      data[48] <= 430227734;
      data[49] <= 506948616;
      data[50] <= 659060556;
      data[51] <= 883997877;
      data[52] <= 958139571;
      data[53] <= 1322822218;
      data[54] <= 1537002063;
      data[55] <= 1747873779;
      data[56] <= 1955562222;
      data[57] <= 2024104815;
      data[58] <= -2067236844;
      data[59] <= -1933114872;
      data[60] <= -1866530822;
      data[61] <= -1538233109;
      data[62] <= -1090935817;
      data[63] <= -965641998;
    end else begin
      if (write_en_i) begin
        data[addr_i] <= wdata_i;
      end
    end
  end
  // Read
  always @(addr_i or clk) begin
    rdata_o = data[addr_i];
  end
endmodule

module axi_master_controller_a4rd32(clk, rst, sram_addr, sram_wdata, sram_wen, sram_rdata, sram_EXCLUSIVE, sram_req, sram_ack, addr, len, start, wen, req, ack, ARADDR, ARVALID, ARREADY, ARLEN, ARSIZE, RVALID, RDATA, RREADY, RLAST, AWADDR, AWVALID, AWREADY, AWLEN, AWSIZE, WVALID, WREADY, WDATA, WLAST, BVALID, BREADY, BRESP);
  input clk;
  input rst;
  output [3:0] sram_addr;
  output [31:0] sram_wdata;
  output sram_wen;
  input [31:0] sram_rdata;
  input sram_EXCLUSIVE;
  output sram_req;
  input sram_ack;
  input [31:0] addr;
  input [3:0] len;
  input [3:0] start;
  input wen;
  input req;
  output ack;
  output [31:0] ARADDR;
  output ARVALID;
  input ARREADY;
  output [7:0] ARLEN;
  output [2:0] ARSIZE;
  input RVALID;
  input [31:0] RDATA;
  output RREADY;
  input RLAST;
  output [31:0] AWADDR;
  output AWVALID;
  input AWREADY;
  output [7:0] AWLEN;
  output [2:0] AWSIZE;
  output WVALID;
  input WREADY;
  output [31:0] WDATA;
  output WLAST;
  input BVALID;
  output BREADY;
  input [1:0] BRESP;
  reg [3:0] sram_addr;
  reg [31:0] sram_wdata;
  reg sram_wen;
  reg sram_req;
  reg ack;
  reg [31:0] ARADDR;
  reg ARVALID;
  reg [7:0] ARLEN;
  reg [2:0] ARSIZE;
  reg RREADY;
  reg [31:0] AWADDR;
  reg AWVALID;
  reg [7:0] AWLEN;
  reg [2:0] AWSIZE;
  reg WVALID;
  reg [31:0] WDATA;
  reg WLAST;
  reg BREADY;

  `define S_IDLE 0
  `define S_ADDR_WAIT 1
  `define S_READ_DATA 2
  `define S_READ_DATA_WAIT 3
  reg [2:0] st;

  reg [4:0] ridx;
  reg read_last;

  always @(posedge clk) begin
    if (rst) begin
      ack <= 0;
      sram_req <= 0;
      sram_wen <= 0;
      st <= `S_IDLE;
      ARADDR <= 0;
      ARVALID <= 0;
      ARLEN <= 0;
      ARSIZE <= 0;
      RREADY <= 0;
      AWADDR <= 0;
      AWVALID <= 0;
      AWLEN <= 0;
      AWSIZE <= 0;
      WVALID <= 0;
      WDATA <= 0;
      WLAST <= 0;
      BREADY <= 0;
    end else begin
      if (sram_EXCLUSIVE) begin
        sram_wen <= (st == `S_READ_DATA && RVALID);
      end
      case (st)
        `S_IDLE: begin
          ack <= 0;
          if (req && !ack) begin
            ridx <= 0;
            st <= `S_ADDR_WAIT;
            ARVALID <= 1;
            ARADDR <= addr;
            ARLEN <= len;
            ARSIZE <= 2;
          end
        end
        `S_ADDR_WAIT: begin
          ack <= 0;
          if (ARREADY) begin
            st <= `S_READ_DATA;
            ARVALID <= 0;
            RREADY <= 1;
          end
        end
        `S_READ_DATA: begin
          if (RVALID) begin
            sram_addr <= start + ridx;
            sram_wdata <= RDATA;
            ridx <= ridx + 1;
            if (sram_EXCLUSIVE) begin
              if (RLAST) begin
                RREADY <= 0;
                ack <= 1;
                st <= `S_IDLE;
              end
            end else begin
              st <= `S_READ_DATA_WAIT;
              sram_req <= 1;
              sram_wen <= 1;
              RREADY <= 0;
              read_last <= RLAST;
            end
          end
        end
        `S_READ_DATA_WAIT: begin
          if (sram_ack) begin
            sram_req <= 0;
            sram_wen <= 0;
            if (read_last) begin
              ack <= 1;
              st <= `S_IDLE;
            end else begin
              st <= `S_READ_DATA;
              RREADY <= 1;
            end
          end
        end
      endcase
    end
  end
endmodule

// Module 1;
module main(clk, rst, buf_ARADDR, buf_ARVALID, buf_ARREADY, buf_ARLEN, buf_ARSIZE, buf_RVALID, buf_RDATA, buf_RREADY, buf_RLAST, buf_AWADDR, buf_AWVALID, buf_AWREADY, buf_AWLEN, buf_AWSIZE, buf_WVALID, buf_WREADY, buf_WDATA, buf_WLAST, buf_BVALID, buf_BREADY, buf_BRESP, sha256_req_valid, sha256_req_ready, sha256_req_busy, sha256_res_valid, sha256_res_ready, sha256_req_0, sha256_req_1, sha256_res_0);
  input clk;
  input rst;
  output [31:0] buf_ARADDR;
  output buf_ARVALID;
  input buf_ARREADY;
  output [7:0] buf_ARLEN;
  output [2:0] buf_ARSIZE;
  input buf_RVALID;
  input [31:0] buf_RDATA;
  output buf_RREADY;
  input buf_RLAST;
  output [31:0] buf_AWADDR;
  output buf_AWVALID;
  input buf_AWREADY;
  output [7:0] buf_AWLEN;
  output [2:0] buf_AWSIZE;
  output buf_WVALID;
  input buf_WREADY;
  output [31:0] buf_WDATA;
  output buf_WLAST;
  input buf_BVALID;
  output buf_BREADY;
  input [1:0] buf_BRESP;
  input sha256_req_valid;
  output sha256_req_ready;
  output sha256_req_busy;
  output sha256_res_valid;
  input sha256_res_ready;
  input [31:0] sha256_req_0;
  input [31:0] sha256_req_1;
  output [255:0] sha256_res_0;
  reg sha256_req_ready;
  reg sha256_req_busy;
  reg sha256_res_valid;
  reg [255:0] sha256_res_0;

  // State decls
  // state names
  `define S_1_1 1
  `define S_1_2 2
  reg [1:0] st_1;

  // state names
  `define S_2_1 1
  `define S_2_6 6
  `define S_2_7 7
  `define S_2_8 8
  `define S_2_9 9
  `define S_2_13 13
  `define S_2_19 19
  `define S_2_20 20
  `define S_2_21 21
  `define S_2_23 23
  `define S_2_26 26
  `define S_2_2 2
  `define S_2_29 29
  `define S_2_33 33
  `define S_2_3 3
  `define S_2_36 36
  `define S_2_37 37
  `define S_2_41 41
  `define S_2_4 4
  `define S_2_44 44
  `define S_2_45 45
  `define S_2_49 49
  `define S_2_5 5
  `define S_2_52 52
  `define S_2_53 53
  `define S_2_57 57
  `define S_2_10 10
  `define S_2_60 60
  `define S_2_61 61
  `define S_2_65 65
  `define S_2_11 11
  `define S_2_68 68
  `define S_2_69 69
  `define S_2_73 73
  `define S_2_12 12
  `define S_2_76 76
  `define S_2_77 77
  `define S_2_81 81
  `define S_2_14 14
  `define S_2_84 84
  `define S_2_85 85
  `define S_2_89 89
  `define S_2_15 15
  `define S_2_92 92
  `define S_2_93 93
  `define S_2_97 97
  `define S_2_16 16
  `define S_2_100 100
  `define S_2_101 101
  `define S_2_105 105
  `define S_2_17 17
  `define S_2_108 108
  `define S_2_109 109
  `define S_2_113 113
  `define S_2_18 18
  `define S_2_116 116
  `define S_2_117 117
  `define S_2_121 121
  `define S_2_22 22
  `define S_2_124 124
  `define S_2_125 125
  `define S_2_129 129
  `define S_2_24 24
  `define S_2_132 132
  `define S_2_133 133
  `define S_2_137 137
  `define S_2_25 25
  `define S_2_140 140
  `define S_2_141 141
  `define S_2_145 145
  `define S_2_27 27
  `define S_2_148 148
  `define S_2_149 149
  `define S_2_153 153
  `define S_2_28 28
  `define S_2_156 156
  `define S_2_157 157
  `define S_2_161 161
  `define S_2_30 30
  `define S_2_164 164
  `define S_2_165 165
  `define S_2_169 169
  `define S_2_31 31
  `define S_2_172 172
  `define S_2_173 173
  `define S_2_177 177
  `define S_2_32 32
  `define S_2_180 180
  `define S_2_181 181
  `define S_2_185 185
  `define S_2_34 34
  `define S_2_188 188
  `define S_2_189 189
  `define S_2_193 193
  `define S_2_35 35
  `define S_2_196 196
  `define S_2_197 197
  `define S_2_201 201
  `define S_2_38 38
  `define S_2_204 204
  `define S_2_205 205
  `define S_2_209 209
  `define S_2_39 39
  `define S_2_212 212
  `define S_2_213 213
  `define S_2_217 217
  `define S_2_40 40
  `define S_2_220 220
  `define S_2_221 221
  `define S_2_225 225
  `define S_2_42 42
  `define S_2_228 228
  `define S_2_229 229
  `define S_2_233 233
  `define S_2_43 43
  `define S_2_236 236
  `define S_2_237 237
  `define S_2_241 241
  `define S_2_46 46
  `define S_2_244 244
  `define S_2_245 245
  `define S_2_249 249
  `define S_2_47 47
  `define S_2_252 252
  `define S_2_253 253
  `define S_2_257 257
  `define S_2_48 48
  `define S_2_260 260
  `define S_2_261 261
  `define S_2_265 265
  `define S_2_50 50
  `define S_2_268 268
  `define S_2_269 269
  `define S_2_273 273
  `define S_2_51 51
  `define S_2_276 276
  `define S_2_277 277
  `define S_2_278 278
  `define S_2_282 282
  `define S_2_288 288
  `define S_2_293 293
  `define S_2_298 298
  `define S_2_303 303
  `define S_2_308 308
  `define S_2_313 313
  `define S_2_318 318
  `define S_2_323 323
  `define S_2_329 329
  `define S_2_330 330
  `define S_2_331 331
  `define S_2_332 332
  `define S_2_333 333
  `define S_2_335 335
  `define S_2_336 336
  `define S_2_339 339
  `define S_2_342 342
  `define S_2_343 343
  `define S_2_346 346
  `define S_2_347 347
  `define S_2_350 350
  `define S_2_351 351
  `define S_2_354 354
  `define S_2_355 355
  `define S_2_357 357
  `define S_2_358 358
  `define S_2_359 359
  `define S_2_360 360
  `define S_2_361 361
  `define S_2_362 362
  `define S_2_364 364
  `define S_2_367 367
  `define S_2_54 54
  `define S_2_368 368
  `define S_2_369 369
  `define S_2_371 371
  `define S_2_374 374
  `define S_2_55 55
  `define S_2_375 375
  `define S_2_378 378
  `define S_2_381 381
  `define S_2_56 56
  `define S_2_382 382
  `define S_2_383 383
  `define S_2_384 384
  `define S_2_386 386
  `define S_2_389 389
  `define S_2_58 58
  `define S_2_390 390
  `define S_2_393 393
  `define S_2_394 394
  `define S_2_396 396
  `define S_2_399 399
  `define S_2_59 59
  `define S_2_400 400
  `define S_2_404 404
  `define S_2_62 62
  `define S_2_405 405
  `define S_2_409 409
  `define S_2_63 63
  `define S_2_410 410
  `define S_2_414 414
  `define S_2_64 64
  `define S_2_415 415
  `define S_2_419 419
  `define S_2_66 66
  `define S_2_420 420
  `define S_2_424 424
  `define S_2_67 67
  `define S_2_425 425
  `define S_2_429 429
  `define S_2_70 70
  `define S_2_430 430
  `define S_2_434 434
  `define S_2_71 71
  `define S_2_435 435
  `define S_2_437 437
  `define S_2_438 438
  `define S_2_439 439
  `define S_2_440 440
  `define S_2_441 441
  `define S_2_442 442
  `define S_2_443 443
  `define S_2_445 445
  `define S_2_446 446
  `define S_2_448 448
  `define S_2_451 451
  `define S_2_72 72
  `define S_2_452 452
  `define S_2_456 456
  `define S_2_460 460
  `define S_2_74 74
  `define S_2_461 461
  `define S_2_465 465
  `define S_2_469 469
  `define S_2_75 75
  `define S_2_470 470
  `define S_2_474 474
  `define S_2_478 478
  `define S_2_78 78
  `define S_2_479 479
  `define S_2_483 483
  `define S_2_487 487
  `define S_2_79 79
  `define S_2_488 488
  `define S_2_492 492
  `define S_2_496 496
  `define S_2_80 80
  `define S_2_497 497
  `define S_2_501 501
  `define S_2_505 505
  `define S_2_82 82
  `define S_2_506 506
  `define S_2_510 510
  `define S_2_514 514
  `define S_2_83 83
  `define S_2_515 515
  `define S_2_519 519
  `define S_2_525 525
  `define S_2_526 526
  `define S_2_528 528
  `define S_2_529 529
  `define S_2_530 530
  `define S_2_532 532
  `define S_2_533 533
  `define S_2_534 534
  `define S_2_542 542
  `define S_2_545 545
  `define S_2_546 546
  `define S_2_547 547
  `define S_2_555 555
  `define S_2_558 558
  `define S_2_559 559
  `define S_2_560 560
  `define S_2_567 567
  `define S_2_568 568
  `define S_2_570 570
  `define S_2_571 571
  `define S_2_572 572
  `define S_2_574 574
  `define S_2_575 575
  `define S_2_576 576
  `define S_2_584 584
  `define S_2_587 587
  `define S_2_588 588
  `define S_2_589 589
  `define S_2_597 597
  `define S_2_600 600
  `define S_2_601 601
  `define S_2_602 602
  `define S_2_609 609
  `define S_2_610 610
  `define S_2_611 611
  `define S_2_613 613
  `define S_2_614 614
  `define S_2_615 615
  `define S_2_618 618
  `define S_2_86 86
  `define S_2_619 619
  `define S_2_622 622
  `define S_2_87 87
  `define S_2_623 623
  `define S_2_624 624
  `define S_2_626 626
  `define S_2_627 627
  `define S_2_629 629
  `define S_2_630 630
  `define S_2_631 631
  `define S_2_632 632
  `define S_2_633 633
  `define S_2_634 634
  `define S_2_635 635
  `define S_2_636 636
  `define S_2_638 638
  `define S_2_639 639
  `define S_2_640 640
  `define S_2_642 642
  `define S_2_643 643
  `define S_2_644 644
  `define S_2_646 646
  `define S_2_649 649
  `define S_2_88 88
  `define S_2_650 650
  `define S_2_652 652
  `define S_2_655 655
  `define S_2_90 90
  `define S_2_656 656
  `define S_2_657 657
  `define S_2_659 659
  `define S_2_660 660
  `define S_2_662 662
  `define S_2_663 663
  `define S_2_664 664
  `define S_2_665 665
  `define S_2_666 666
  `define S_2_667 667
  `define S_2_668 668
  `define S_2_669 669
  `define S_2_671 671
  `define S_2_672 672
  `define S_2_673 673
  `define S_2_675 675
  `define S_2_676 676
  `define S_2_677 677
  `define S_2_679 679
  `define S_2_682 682
  `define S_2_91 91
  `define S_2_683 683
  `define S_2_685 685
  `define S_2_688 688
  `define S_2_94 94
  `define S_2_689 689
  `define S_2_690 690
  `define S_2_692 692
  `define S_2_693 693
  `define S_2_695 695
  `define S_2_696 696
  `define S_2_697 697
  `define S_2_698 698
  `define S_2_699 699
  `define S_2_700 700
  `define S_2_701 701
  `define S_2_702 702
  `define S_2_704 704
  `define S_2_705 705
  `define S_2_706 706
  `define S_2_708 708
  `define S_2_709 709
  `define S_2_710 710
  `define S_2_712 712
  `define S_2_715 715
  `define S_2_95 95
  `define S_2_716 716
  `define S_2_718 718
  `define S_2_721 721
  `define S_2_96 96
  `define S_2_722 722
  `define S_2_723 723
  `define S_2_725 725
  `define S_2_726 726
  `define S_2_728 728
  `define S_2_729 729
  `define S_2_730 730
  `define S_2_731 731
  `define S_2_732 732
  `define S_2_733 733
  `define S_2_734 734
  `define S_2_735 735
  `define S_2_737 737
  `define S_2_738 738
  `define S_2_739 739
  `define S_2_741 741
  `define S_2_742 742
  `define S_2_743 743
  `define S_2_745 745
  `define S_2_748 748
  `define S_2_98 98
  `define S_2_749 749
  `define S_2_751 751
  `define S_2_754 754
  `define S_2_99 99
  `define S_2_755 755
  `define S_2_756 756
  `define S_2_758 758
  `define S_2_759 759
  `define S_2_761 761
  `define S_2_762 762
  `define S_2_763 763
  `define S_2_764 764
  `define S_2_765 765
  `define S_2_766 766
  `define S_2_767 767
  `define S_2_768 768
  `define S_2_770 770
  `define S_2_771 771
  `define S_2_772 772
  `define S_2_774 774
  `define S_2_775 775
  `define S_2_776 776
  `define S_2_778 778
  `define S_2_781 781
  `define S_2_102 102
  `define S_2_782 782
  `define S_2_784 784
  `define S_2_787 787
  `define S_2_103 103
  `define S_2_788 788
  `define S_2_789 789
  `define S_2_791 791
  `define S_2_792 792
  `define S_2_794 794
  `define S_2_795 795
  `define S_2_796 796
  `define S_2_797 797
  `define S_2_798 798
  `define S_2_799 799
  `define S_2_800 800
  `define S_2_801 801
  `define S_2_803 803
  `define S_2_804 804
  `define S_2_805 805
  `define S_2_807 807
  `define S_2_808 808
  `define S_2_809 809
  `define S_2_811 811
  `define S_2_814 814
  `define S_2_104 104
  `define S_2_815 815
  `define S_2_817 817
  `define S_2_820 820
  `define S_2_106 106
  `define S_2_821 821
  `define S_2_822 822
  `define S_2_824 824
  `define S_2_825 825
  `define S_2_827 827
  `define S_2_828 828
  `define S_2_829 829
  `define S_2_830 830
  `define S_2_831 831
  `define S_2_832 832
  `define S_2_833 833
  `define S_2_834 834
  `define S_2_836 836
  `define S_2_837 837
  `define S_2_838 838
  `define S_2_840 840
  `define S_2_841 841
  `define S_2_842 842
  `define S_2_844 844
  `define S_2_847 847
  `define S_2_107 107
  `define S_2_848 848
  `define S_2_850 850
  `define S_2_853 853
  `define S_2_110 110
  `define S_2_854 854
  `define S_2_855 855
  `define S_2_857 857
  `define S_2_858 858
  `define S_2_860 860
  `define S_2_861 861
  `define S_2_862 862
  `define S_2_863 863
  `define S_2_864 864
  `define S_2_865 865
  `define S_2_866 866
  `define S_2_867 867
  `define S_2_868 868
  `define S_2_869 869
  `define S_2_870 870
  `define S_2_871 871
  `define S_2_872 872
  `define S_2_873 873
  `define S_2_874 874
  `define S_2_875 875
  `define S_2_882 882
  `define S_2_883 883
  `define S_2_885 885
  `define S_2_886 886
  `define S_2_887 887
  `define S_2_889 889
  `define S_2_890 890
  `define S_2_891 891
  `define S_2_892 892
  `define S_2_900 900
  `define S_2_903 903
  `define S_2_904 904
  `define S_2_905 905
  `define S_2_913 913
  `define S_2_916 916
  `define S_2_917 917
  `define S_2_918 918
  `define S_2_926 926
  `define S_2_929 929
  `define S_2_930 930
  `define S_2_931 931
  `define S_2_937 937
  `define S_2_938 938
  `define S_2_939 939
  `define S_2_940 940
  `define S_2_947 947
  `define S_2_948 948
  `define S_2_950 950
  `define S_2_951 951
  `define S_2_952 952
  `define S_2_954 954
  `define S_2_955 955
  `define S_2_956 956
  `define S_2_957 957
  `define S_2_965 965
  `define S_2_968 968
  `define S_2_969 969
  `define S_2_970 970
  `define S_2_978 978
  `define S_2_981 981
  `define S_2_982 982
  `define S_2_983 983
  `define S_2_991 991
  `define S_2_994 994
  `define S_2_995 995
  `define S_2_996 996
  `define S_2_1002 1002
  `define S_2_1003 1003
  `define S_2_1004 1004
  `define S_2_1005 1005
  `define S_2_1006 1006
  `define S_2_1013 1013
  `define S_2_1014 1014
  `define S_2_1016 1016
  `define S_2_1017 1017
  `define S_2_1018 1018
  `define S_2_1020 1020
  `define S_2_1021 1021
  `define S_2_1022 1022
  `define S_2_1023 1023
  `define S_2_1031 1031
  `define S_2_1034 1034
  `define S_2_1035 1035
  `define S_2_1036 1036
  `define S_2_1044 1044
  `define S_2_1047 1047
  `define S_2_1048 1048
  `define S_2_1049 1049
  `define S_2_1057 1057
  `define S_2_1060 1060
  `define S_2_1061 1061
  `define S_2_1062 1062
  `define S_2_1068 1068
  `define S_2_1069 1069
  `define S_2_1070 1070
  `define S_2_1071 1071
  `define S_2_1078 1078
  `define S_2_1079 1079
  `define S_2_1081 1081
  `define S_2_1082 1082
  `define S_2_1083 1083
  `define S_2_1085 1085
  `define S_2_1086 1086
  `define S_2_1087 1087
  `define S_2_1088 1088
  `define S_2_1096 1096
  `define S_2_1099 1099
  `define S_2_1100 1100
  `define S_2_1101 1101
  `define S_2_1109 1109
  `define S_2_1112 1112
  `define S_2_1113 1113
  `define S_2_1114 1114
  `define S_2_1122 1122
  `define S_2_1125 1125
  `define S_2_1126 1126
  `define S_2_1127 1127
  `define S_2_1133 1133
  `define S_2_1134 1134
  `define S_2_1135 1135
  `define S_2_1136 1136
  `define S_2_1137 1137
  `define S_2_1144 1144
  `define S_2_1145 1145
  `define S_2_1147 1147
  `define S_2_1148 1148
  `define S_2_1149 1149
  `define S_2_1151 1151
  `define S_2_1152 1152
  `define S_2_1153 1153
  `define S_2_1154 1154
  `define S_2_1162 1162
  `define S_2_1165 1165
  `define S_2_1166 1166
  `define S_2_1167 1167
  `define S_2_1175 1175
  `define S_2_1178 1178
  `define S_2_1179 1179
  `define S_2_1180 1180
  `define S_2_1188 1188
  `define S_2_1191 1191
  `define S_2_1192 1192
  `define S_2_1193 1193
  `define S_2_1199 1199
  `define S_2_1200 1200
  `define S_2_1201 1201
  `define S_2_1202 1202
  `define S_2_1209 1209
  `define S_2_1210 1210
  `define S_2_1212 1212
  `define S_2_1213 1213
  `define S_2_1214 1214
  `define S_2_1216 1216
  `define S_2_1217 1217
  `define S_2_1218 1218
  `define S_2_1219 1219
  `define S_2_1227 1227
  `define S_2_1230 1230
  `define S_2_1231 1231
  `define S_2_1232 1232
  `define S_2_1240 1240
  `define S_2_1243 1243
  `define S_2_1244 1244
  `define S_2_1245 1245
  `define S_2_1253 1253
  `define S_2_1256 1256
  `define S_2_1257 1257
  `define S_2_1258 1258
  `define S_2_1264 1264
  `define S_2_1265 1265
  `define S_2_1266 1266
  `define S_2_1267 1267
  `define S_2_1268 1268
  `define S_2_1275 1275
  `define S_2_1276 1276
  `define S_2_1278 1278
  `define S_2_1279 1279
  `define S_2_1280 1280
  `define S_2_1282 1282
  `define S_2_1283 1283
  `define S_2_1284 1284
  `define S_2_1285 1285
  `define S_2_1293 1293
  `define S_2_1296 1296
  `define S_2_1297 1297
  `define S_2_1298 1298
  `define S_2_1306 1306
  `define S_2_1309 1309
  `define S_2_1310 1310
  `define S_2_1311 1311
  `define S_2_1319 1319
  `define S_2_1322 1322
  `define S_2_1323 1323
  `define S_2_1324 1324
  `define S_2_1330 1330
  `define S_2_1331 1331
  `define S_2_1332 1332
  `define S_2_1333 1333
  `define S_2_1340 1340
  `define S_2_1341 1341
  `define S_2_1343 1343
  `define S_2_1344 1344
  `define S_2_1345 1345
  `define S_2_1347 1347
  `define S_2_1348 1348
  `define S_2_1349 1349
  `define S_2_1350 1350
  `define S_2_1358 1358
  `define S_2_1361 1361
  `define S_2_1362 1362
  `define S_2_1363 1363
  `define S_2_1371 1371
  `define S_2_1374 1374
  `define S_2_1375 1375
  `define S_2_1376 1376
  `define S_2_1384 1384
  `define S_2_1387 1387
  `define S_2_1388 1388
  `define S_2_1389 1389
  `define S_2_1395 1395
  `define S_2_1396 1396
  `define S_2_1397 1397
  `define S_2_1398 1398
  `define S_2_1399 1399
  `define S_2_1406 1406
  `define S_2_1407 1407
  `define S_2_1409 1409
  `define S_2_1410 1410
  `define S_2_1411 1411
  `define S_2_1413 1413
  `define S_2_1414 1414
  `define S_2_1415 1415
  `define S_2_1416 1416
  `define S_2_1424 1424
  `define S_2_1427 1427
  `define S_2_1428 1428
  `define S_2_1429 1429
  `define S_2_1437 1437
  `define S_2_1440 1440
  `define S_2_1441 1441
  `define S_2_1442 1442
  `define S_2_1450 1450
  `define S_2_1453 1453
  `define S_2_1454 1454
  `define S_2_1455 1455
  `define S_2_1461 1461
  `define S_2_1462 1462
  `define S_2_1463 1463
  `define S_2_1464 1464
  `define S_2_1471 1471
  `define S_2_1472 1472
  `define S_2_1474 1474
  `define S_2_1475 1475
  `define S_2_1476 1476
  `define S_2_1478 1478
  `define S_2_1479 1479
  `define S_2_1480 1480
  `define S_2_1481 1481
  `define S_2_1489 1489
  `define S_2_1492 1492
  `define S_2_1493 1493
  `define S_2_1494 1494
  `define S_2_1502 1502
  `define S_2_1505 1505
  `define S_2_1506 1506
  `define S_2_1507 1507
  `define S_2_1515 1515
  `define S_2_1518 1518
  `define S_2_1519 1519
  `define S_2_1520 1520
  `define S_2_1526 1526
  `define S_2_1527 1527
  `define S_2_1528 1528
  `define S_2_1529 1529
  `define S_2_1530 1530
  `define S_2_1537 1537
  `define S_2_1538 1538
  `define S_2_1540 1540
  `define S_2_1541 1541
  `define S_2_1542 1542
  `define S_2_1544 1544
  `define S_2_1545 1545
  `define S_2_1546 1546
  `define S_2_1547 1547
  `define S_2_1555 1555
  `define S_2_1558 1558
  `define S_2_1559 1559
  `define S_2_1560 1560
  `define S_2_1568 1568
  `define S_2_1571 1571
  `define S_2_1572 1572
  `define S_2_1573 1573
  `define S_2_1581 1581
  `define S_2_1584 1584
  `define S_2_1585 1585
  `define S_2_1586 1586
  `define S_2_1592 1592
  `define S_2_1593 1593
  `define S_2_1594 1594
  `define S_2_1595 1595
  `define S_2_1602 1602
  `define S_2_1603 1603
  `define S_2_1605 1605
  `define S_2_1606 1606
  `define S_2_1607 1607
  `define S_2_1609 1609
  `define S_2_1610 1610
  `define S_2_1611 1611
  `define S_2_1612 1612
  `define S_2_1620 1620
  `define S_2_1623 1623
  `define S_2_1624 1624
  `define S_2_1625 1625
  `define S_2_1633 1633
  `define S_2_1636 1636
  `define S_2_1637 1637
  `define S_2_1638 1638
  `define S_2_1646 1646
  `define S_2_1649 1649
  `define S_2_1650 1650
  `define S_2_1651 1651
  `define S_2_1657 1657
  `define S_2_1658 1658
  `define S_2_1659 1659
  `define S_2_1660 1660
  `define S_2_1661 1661
  `define S_2_1668 1668
  `define S_2_1669 1669
  `define S_2_1671 1671
  `define S_2_1672 1672
  `define S_2_1673 1673
  `define S_2_1675 1675
  `define S_2_1676 1676
  `define S_2_1677 1677
  `define S_2_1678 1678
  `define S_2_1686 1686
  `define S_2_1689 1689
  `define S_2_1690 1690
  `define S_2_1691 1691
  `define S_2_1699 1699
  `define S_2_1702 1702
  `define S_2_1703 1703
  `define S_2_1704 1704
  `define S_2_1712 1712
  `define S_2_1715 1715
  `define S_2_1716 1716
  `define S_2_1717 1717
  `define S_2_1723 1723
  `define S_2_1724 1724
  `define S_2_1725 1725
  `define S_2_1726 1726
  `define S_2_1733 1733
  `define S_2_1734 1734
  `define S_2_1736 1736
  `define S_2_1737 1737
  `define S_2_1738 1738
  `define S_2_1740 1740
  `define S_2_1741 1741
  `define S_2_1742 1742
  `define S_2_1743 1743
  `define S_2_1751 1751
  `define S_2_1754 1754
  `define S_2_1755 1755
  `define S_2_1756 1756
  `define S_2_1764 1764
  `define S_2_1767 1767
  `define S_2_1768 1768
  `define S_2_1769 1769
  `define S_2_1777 1777
  `define S_2_1780 1780
  `define S_2_1781 1781
  `define S_2_1782 1782
  `define S_2_1788 1788
  `define S_2_1789 1789
  `define S_2_1790 1790
  `define S_2_1791 1791
  `define S_2_1792 1792
  `define S_2_1799 1799
  `define S_2_1800 1800
  `define S_2_1802 1802
  `define S_2_1803 1803
  `define S_2_1804 1804
  `define S_2_1806 1806
  `define S_2_1807 1807
  `define S_2_1808 1808
  `define S_2_1809 1809
  `define S_2_1817 1817
  `define S_2_1820 1820
  `define S_2_1821 1821
  `define S_2_1822 1822
  `define S_2_1830 1830
  `define S_2_1833 1833
  `define S_2_1834 1834
  `define S_2_1835 1835
  `define S_2_1843 1843
  `define S_2_1846 1846
  `define S_2_1847 1847
  `define S_2_1848 1848
  `define S_2_1854 1854
  `define S_2_1855 1855
  `define S_2_1856 1856
  `define S_2_1857 1857
  `define S_2_1864 1864
  `define S_2_1865 1865
  `define S_2_1867 1867
  `define S_2_1868 1868
  `define S_2_1869 1869
  `define S_2_1871 1871
  `define S_2_1872 1872
  `define S_2_1873 1873
  `define S_2_1874 1874
  `define S_2_1882 1882
  `define S_2_1885 1885
  `define S_2_1886 1886
  `define S_2_1887 1887
  `define S_2_1895 1895
  `define S_2_1898 1898
  `define S_2_1899 1899
  `define S_2_1900 1900
  `define S_2_1908 1908
  `define S_2_1911 1911
  `define S_2_1912 1912
  `define S_2_1913 1913
  `define S_2_1919 1919
  `define S_2_1920 1920
  `define S_2_1921 1921
  `define S_2_1922 1922
  `define S_2_1923 1923
  `define S_2_task_idle 1924
  reg [11:0] st_2;

  // State vars
  // Registers
  reg  [31:0] r__29_493;
  reg  [31:0] arg_177_561;
  reg  [31:0] r1_ror32_17_178_565;
  reg  [16:0] r3_ror32_17_179_562;
  reg  [14:0] r6_ror32_17_180_563;
  reg  [31:0] r2_ror32_17_181_564;
  reg  [12:0] r6_ror32_19_190_568;
  reg  [31:0] arg_187_566;
  reg  [31:0] r1_ror32_19_188_570;
  reg  [18:0] r3_ror32_19_189_567;
  reg  [31:0] r2_ror32_19_191_569;
  reg  [31:0] x_224_554;
  reg  [31:0] r1_s1_225_560;
  reg  [31:0] r4_s1_226_555;
  reg  [31:0] r6_s1_227_556;
  reg  [31:0] r3_s1_228_557;
  reg  [31:0] r8_s1_229_558;
  reg  [31:0] r2_s1_230_559;
  reg  [31:0] arg_212_578;
  reg  [31:0] r1_ror32_7_213_582;
  reg  [6:0] r3_ror32_7_214_579;
  reg  [24:0] r6_ror32_7_215_580;
  reg  [31:0] r2_ror32_7_216_581;
  reg  [31:0] arg_182_583;
  reg  [31:0] r1_ror32_18_183_587;
  reg  [17:0] r3_ror32_18_184_584;
  reg  [13:0] r6_ror32_18_185_585;
  reg  [31:0] r2_ror32_18_186_586;
  reg  [31:0] r8_s0_222_575;
  reg  [31:0] r2_s0_223_576;
  reg  [31:0] x_217_571;
  reg  [31:0] r1_s0_218_577;
  reg  [31:0] r4_s0_219_572;
  reg  [31:0] r6_s0_220_573;
  reg  [31:0] r3_s0_221_574;
  reg  [31:0] arg_207_732;
  reg  [31:0] r1_ror32_6_208_736;
  reg  [5:0] r3_ror32_6_209_733;
  reg  [25:0] r6_ror32_6_210_734;
  reg  [31:0] r2_ror32_6_211_735;
  reg  [31:0] arg_167_737;
  reg  [31:0] r1_ror32_11_168_741;
  reg  [10:0] r3_ror32_11_169_738;
  reg  [20:0] r6_ror32_11_170_739;
  reg  [31:0] r2_ror32_11_171_740;
  reg  [31:0] arg_202_742;
  reg  [31:0] r1_ror32_25_203_746;
  reg  [24:0] r3_ror32_25_204_743;
  reg  [6:0] r6_ror32_25_205_744;
  reg  [31:0] r2_ror32_25_206_745;
  reg  [31:0] x_22_725;
  reg  [31:0] r1_e1_23_731;
  reg  [31:0] r4_e1_24_726;
  reg  [31:0] r6_e1_25_727;
  reg  [31:0] r3_e1_26_728;
  reg  [31:0] r8_e1_27_729;
  reg  [31:0] r2_e1_28_730;
  reg  [31:0] x_0_750;
  reg  [31:0] y_1_747;
  reg  [31:0] z_2_748;
  reg  [31:0] r3_Ch_3_753;
  reg  [31:0] r6_Ch_4_749;
  reg  [31:0] r5_Ch_5_751;
  reg  [31:0] r4_Ch_6_752;
  reg  [31:0] arg_192_761;
  reg  [31:0] r1_ror32_2_193_765;
  reg  [1:0] r3_ror32_2_194_762;
  reg  [29:0] r6_ror32_2_195_763;
  reg  [31:0] r2_ror32_2_196_764;
  reg  [31:0] arg_172_766;
  reg  [31:0] r1_ror32_13_173_770;
  reg  [12:0] r3_ror32_13_174_767;
  reg  [18:0] r6_ror32_13_175_768;
  reg  [31:0] r2_ror32_13_176_769;
  reg  [31:0] arg_197_771;
  reg  [31:0] r1_ror32_22_198_775;
  reg  [21:0] r3_ror32_22_199_772;
  reg  [9:0] r6_ror32_22_200_773;
  reg  [31:0] r2_ror32_22_201_774;
  reg  [31:0] x_15_754;
  reg  [31:0] r1_e0_16_760;
  reg  [31:0] r4_e0_17_755;
  reg  [31:0] r6_e0_18_756;
  reg  [31:0] r3_e0_19_757;
  reg  [31:0] r8_e0_20_758;
  reg  [31:0] r2_e0_21_759;
  reg  [31:0] x_7_776;
  reg  [31:0] y_8_777;
  reg  [31:0] z_9_780;
  reg  [31:0] r3_Maj_10_783;
  reg  [31:0] r5_Maj_11_778;
  reg  [31:0] r7_Maj_12_779;
  reg  [31:0] r6_Maj_13_781;
  reg  [31:0] r4_Maj_14_782;
  reg  [31:0] arg_207_791;
  reg  [31:0] r1_ror32_6_208_795;
  reg  [5:0] r3_ror32_6_209_792;
  reg  [25:0] r6_ror32_6_210_793;
  reg  [31:0] r2_ror32_6_211_794;
  reg  [31:0] arg_167_796;
  reg  [31:0] r1_ror32_11_168_800;
  reg  [10:0] r3_ror32_11_169_797;
  reg  [20:0] r6_ror32_11_170_798;
  reg  [31:0] r2_ror32_11_171_799;
  reg  [31:0] arg_202_801;
  reg  [31:0] r1_ror32_25_203_805;
  reg  [24:0] r3_ror32_25_204_802;
  reg  [6:0] r6_ror32_25_205_803;
  reg  [31:0] r2_ror32_25_206_804;
  reg  [31:0] x_22_784;
  reg  [31:0] r1_e1_23_790;
  reg  [31:0] r4_e1_24_785;
  reg  [31:0] r6_e1_25_786;
  reg  [31:0] r3_e1_26_787;
  reg  [31:0] r8_e1_27_788;
  reg  [31:0] r2_e1_28_789;
  reg  [31:0] x_0_809;
  reg  [31:0] y_1_806;
  reg  [31:0] z_2_807;
  reg  [31:0] r3_Ch_3_812;
  reg  [31:0] r6_Ch_4_808;
  reg  [31:0] r5_Ch_5_810;
  reg  [31:0] r4_Ch_6_811;
  reg  [31:0] arg_192_820;
  reg  [31:0] r1_ror32_2_193_824;
  reg  [1:0] r3_ror32_2_194_821;
  reg  [29:0] r6_ror32_2_195_822;
  reg  [31:0] r2_ror32_2_196_823;
  reg  [31:0] arg_172_825;
  reg  [31:0] r1_ror32_13_173_829;
  reg  [12:0] r3_ror32_13_174_826;
  reg  [18:0] r6_ror32_13_175_827;
  reg  [31:0] r2_ror32_13_176_828;
  reg  [31:0] arg_197_830;
  reg  [31:0] r1_ror32_22_198_834;
  reg  [21:0] r3_ror32_22_199_831;
  reg  [9:0] r6_ror32_22_200_832;
  reg  [31:0] r2_ror32_22_201_833;
  reg  [31:0] x_15_813;
  reg  [31:0] r1_e0_16_819;
  reg  [31:0] r4_e0_17_814;
  reg  [31:0] r6_e0_18_815;
  reg  [31:0] r3_e0_19_816;
  reg  [31:0] r8_e0_20_817;
  reg  [31:0] r2_e0_21_818;
  reg  [31:0] x_7_835;
  reg  [31:0] y_8_836;
  reg  [31:0] z_9_839;
  reg  [31:0] r3_Maj_10_842;
  reg  [31:0] r5_Maj_11_837;
  reg  [31:0] r7_Maj_12_838;
  reg  [31:0] r6_Maj_13_840;
  reg  [31:0] r4_Maj_14_841;
  reg  [31:0] arg_207_850;
  reg  [31:0] r1_ror32_6_208_854;
  reg  [5:0] r3_ror32_6_209_851;
  reg  [25:0] r6_ror32_6_210_852;
  reg  [31:0] r2_ror32_6_211_853;
  reg  [31:0] arg_167_855;
  reg  [31:0] r1_ror32_11_168_859;
  reg  [10:0] r3_ror32_11_169_856;
  reg  [20:0] r6_ror32_11_170_857;
  reg  [31:0] r2_ror32_11_171_858;
  reg  [31:0] arg_202_860;
  reg  [31:0] r1_ror32_25_203_864;
  reg  [24:0] r3_ror32_25_204_861;
  reg  [6:0] r6_ror32_25_205_862;
  reg  [31:0] r2_ror32_25_206_863;
  reg  [31:0] x_22_843;
  reg  [31:0] r1_e1_23_849;
  reg  [31:0] r4_e1_24_844;
  reg  [31:0] r6_e1_25_845;
  reg  [31:0] r3_e1_26_846;
  reg  [31:0] r8_e1_27_847;
  reg  [31:0] r2_e1_28_848;
  reg  [31:0] x_0_868;
  reg  [31:0] y_1_865;
  reg  [31:0] z_2_866;
  reg  [31:0] r3_Ch_3_871;
  reg  [31:0] r6_Ch_4_867;
  reg  [31:0] r5_Ch_5_869;
  reg  [31:0] r4_Ch_6_870;
  reg  [31:0] arg_192_879;
  reg  [31:0] r1_ror32_2_193_883;
  reg  [1:0] r3_ror32_2_194_880;
  reg  [29:0] r6_ror32_2_195_881;
  reg  [31:0] r2_ror32_2_196_882;
  reg  [31:0] arg_172_884;
  reg  [31:0] r1_ror32_13_173_888;
  reg  [12:0] r3_ror32_13_174_885;
  reg  [18:0] r6_ror32_13_175_886;
  reg  [31:0] r2_ror32_13_176_887;
  reg  [31:0] arg_197_889;
  reg  [31:0] r1_ror32_22_198_893;
  reg  [21:0] r3_ror32_22_199_890;
  reg  [9:0] r6_ror32_22_200_891;
  reg  [31:0] r2_ror32_22_201_892;
  reg  [31:0] x_15_872;
  reg  [31:0] r1_e0_16_878;
  reg  [31:0] r4_e0_17_873;
  reg  [31:0] r6_e0_18_874;
  reg  [31:0] r3_e0_19_875;
  reg  [31:0] r8_e0_20_876;
  reg  [31:0] r2_e0_21_877;
  reg  [31:0] x_7_894;
  reg  [31:0] y_8_895;
  reg  [31:0] z_9_898;
  reg  [31:0] r3_Maj_10_901;
  reg  [31:0] r5_Maj_11_896;
  reg  [31:0] r7_Maj_12_897;
  reg  [31:0] r6_Maj_13_899;
  reg  [31:0] r4_Maj_14_900;
  reg  [31:0] arg_207_909;
  reg  [31:0] r1_ror32_6_208_913;
  reg  [5:0] r3_ror32_6_209_910;
  reg  [25:0] r6_ror32_6_210_911;
  reg  [31:0] r2_ror32_6_211_912;
  reg  [31:0] arg_167_914;
  reg  [31:0] r1_ror32_11_168_918;
  reg  [10:0] r3_ror32_11_169_915;
  reg  [20:0] r6_ror32_11_170_916;
  reg  [31:0] r2_ror32_11_171_917;
  reg  [31:0] arg_202_919;
  reg  [31:0] r1_ror32_25_203_923;
  reg  [24:0] r3_ror32_25_204_920;
  reg  [6:0] r6_ror32_25_205_921;
  reg  [31:0] r2_ror32_25_206_922;
  reg  [31:0] x_22_902;
  reg  [31:0] r1_e1_23_908;
  reg  [31:0] r4_e1_24_903;
  reg  [31:0] r6_e1_25_904;
  reg  [31:0] r3_e1_26_905;
  reg  [31:0] r8_e1_27_906;
  reg  [31:0] r2_e1_28_907;
  reg  [31:0] x_0_927;
  reg  [31:0] y_1_924;
  reg  [31:0] z_2_925;
  reg  [31:0] r3_Ch_3_930;
  reg  [31:0] r6_Ch_4_926;
  reg  [31:0] r5_Ch_5_928;
  reg  [31:0] r4_Ch_6_929;
  reg  [31:0] arg_192_938;
  reg  [31:0] r1_ror32_2_193_942;
  reg  [1:0] r3_ror32_2_194_939;
  reg  [29:0] r6_ror32_2_195_940;
  reg  [31:0] r2_ror32_2_196_941;
  reg  [31:0] arg_172_943;
  reg  [31:0] r1_ror32_13_173_947;
  reg  [12:0] r3_ror32_13_174_944;
  reg  [18:0] r6_ror32_13_175_945;
  reg  [31:0] r2_ror32_13_176_946;
  reg  [31:0] arg_197_948;
  reg  [31:0] r1_ror32_22_198_952;
  reg  [21:0] r3_ror32_22_199_949;
  reg  [9:0] r6_ror32_22_200_950;
  reg  [31:0] r2_ror32_22_201_951;
  reg  [31:0] x_15_931;
  reg  [31:0] r1_e0_16_937;
  reg  [31:0] r4_e0_17_932;
  reg  [31:0] r6_e0_18_933;
  reg  [31:0] r3_e0_19_934;
  reg  [31:0] r8_e0_20_935;
  reg  [31:0] r2_e0_21_936;
  reg  [31:0] x_7_953;
  reg  [31:0] y_8_954;
  reg  [31:0] z_9_957;
  reg  [31:0] r3_Maj_10_960;
  reg  [31:0] r5_Maj_11_955;
  reg  [31:0] r7_Maj_12_956;
  reg  [31:0] r6_Maj_13_958;
  reg  [31:0] r4_Maj_14_959;
  reg  [31:0] arg_207_968;
  reg  [31:0] r1_ror32_6_208_972;
  reg  [5:0] r3_ror32_6_209_969;
  reg  [25:0] r6_ror32_6_210_970;
  reg  [31:0] r2_ror32_6_211_971;
  reg  [31:0] arg_167_973;
  reg  [31:0] r1_ror32_11_168_977;
  reg  [10:0] r3_ror32_11_169_974;
  reg  [20:0] r6_ror32_11_170_975;
  reg  [31:0] r2_ror32_11_171_976;
  reg  [31:0] arg_202_978;
  reg  [31:0] r1_ror32_25_203_982;
  reg  [24:0] r3_ror32_25_204_979;
  reg  [6:0] r6_ror32_25_205_980;
  reg  [31:0] r2_ror32_25_206_981;
  reg  [31:0] x_22_961;
  reg  [31:0] r1_e1_23_967;
  reg  [31:0] r4_e1_24_962;
  reg  [31:0] r6_e1_25_963;
  reg  [31:0] r3_e1_26_964;
  reg  [31:0] r8_e1_27_965;
  reg  [31:0] r2_e1_28_966;
  reg  [31:0] x_0_986;
  reg  [31:0] y_1_983;
  reg  [31:0] z_2_984;
  reg  [31:0] r3_Ch_3_989;
  reg  [31:0] r6_Ch_4_985;
  reg  [31:0] r5_Ch_5_987;
  reg  [31:0] r4_Ch_6_988;
  reg  [31:0] arg_192_997;
  reg  [31:0] r1_ror32_2_193_1001;
  reg  [1:0] r3_ror32_2_194_998;
  reg  [29:0] r6_ror32_2_195_999;
  reg  [31:0] r2_ror32_2_196_1000;
  reg  [31:0] arg_172_1002;
  reg  [31:0] r1_ror32_13_173_1006;
  reg  [12:0] r3_ror32_13_174_1003;
  reg  [18:0] r6_ror32_13_175_1004;
  reg  [31:0] r2_ror32_13_176_1005;
  reg  [31:0] arg_197_1007;
  reg  [31:0] r1_ror32_22_198_1011;
  reg  [21:0] r3_ror32_22_199_1008;
  reg  [9:0] r6_ror32_22_200_1009;
  reg  [31:0] r2_ror32_22_201_1010;
  reg  [31:0] x_15_990;
  reg  [31:0] r1_e0_16_996;
  reg  [31:0] r4_e0_17_991;
  reg  [31:0] r6_e0_18_992;
  reg  [31:0] r3_e0_19_993;
  reg  [31:0] r8_e0_20_994;
  reg  [31:0] r2_e0_21_995;
  reg  [31:0] x_7_1012;
  reg  [31:0] y_8_1013;
  reg  [31:0] z_9_1016;
  reg  [31:0] r3_Maj_10_1019;
  reg  [31:0] r5_Maj_11_1014;
  reg  [31:0] r7_Maj_12_1015;
  reg  [31:0] r6_Maj_13_1017;
  reg  [31:0] r4_Maj_14_1018;
  reg  [31:0] arg_207_1027;
  reg  [31:0] r1_ror32_6_208_1031;
  reg  [5:0] r3_ror32_6_209_1028;
  reg  [25:0] r6_ror32_6_210_1029;
  reg  [31:0] r2_ror32_6_211_1030;
  reg  [31:0] arg_167_1032;
  reg  [31:0] r1_ror32_11_168_1036;
  reg  [10:0] r3_ror32_11_169_1033;
  reg  [20:0] r6_ror32_11_170_1034;
  reg  [31:0] r2_ror32_11_171_1035;
  reg  [31:0] arg_202_1037;
  reg  [31:0] r1_ror32_25_203_1041;
  reg  [24:0] r3_ror32_25_204_1038;
  reg  [6:0] r6_ror32_25_205_1039;
  reg  [31:0] r2_ror32_25_206_1040;
  reg  [31:0] x_22_1020;
  reg  [31:0] r1_e1_23_1026;
  reg  [31:0] r4_e1_24_1021;
  reg  [31:0] r6_e1_25_1022;
  reg  [31:0] r3_e1_26_1023;
  reg  [31:0] r8_e1_27_1024;
  reg  [31:0] r2_e1_28_1025;
  reg  [31:0] x_0_1045;
  reg  [31:0] y_1_1042;
  reg  [31:0] z_2_1043;
  reg  [31:0] r3_Ch_3_1048;
  reg  [31:0] r6_Ch_4_1044;
  reg  [31:0] r5_Ch_5_1046;
  reg  [31:0] r4_Ch_6_1047;
  reg  [31:0] arg_192_1056;
  reg  [31:0] r1_ror32_2_193_1060;
  reg  [1:0] r3_ror32_2_194_1057;
  reg  [29:0] r6_ror32_2_195_1058;
  reg  [31:0] r2_ror32_2_196_1059;
  reg  [31:0] arg_172_1061;
  reg  [31:0] r1_ror32_13_173_1065;
  reg  [12:0] r3_ror32_13_174_1062;
  reg  [18:0] r6_ror32_13_175_1063;
  reg  [31:0] r2_ror32_13_176_1064;
  reg  [31:0] arg_197_1066;
  reg  [31:0] r1_ror32_22_198_1070;
  reg  [21:0] r3_ror32_22_199_1067;
  reg  [9:0] r6_ror32_22_200_1068;
  reg  [31:0] r2_ror32_22_201_1069;
  reg  [31:0] x_15_1049;
  reg  [31:0] r1_e0_16_1055;
  reg  [31:0] r4_e0_17_1050;
  reg  [31:0] r6_e0_18_1051;
  reg  [31:0] r3_e0_19_1052;
  reg  [31:0] r8_e0_20_1053;
  reg  [31:0] r2_e0_21_1054;
  reg  [31:0] x_7_1071;
  reg  [31:0] y_8_1072;
  reg  [31:0] z_9_1075;
  reg  [31:0] r3_Maj_10_1078;
  reg  [31:0] r5_Maj_11_1073;
  reg  [31:0] r7_Maj_12_1074;
  reg  [31:0] r6_Maj_13_1076;
  reg  [31:0] r4_Maj_14_1077;
  reg  [31:0] arg_207_1086;
  reg  [31:0] r1_ror32_6_208_1090;
  reg  [5:0] r3_ror32_6_209_1087;
  reg  [25:0] r6_ror32_6_210_1088;
  reg  [31:0] r2_ror32_6_211_1089;
  reg  [31:0] arg_167_1091;
  reg  [31:0] r1_ror32_11_168_1095;
  reg  [10:0] r3_ror32_11_169_1092;
  reg  [20:0] r6_ror32_11_170_1093;
  reg  [31:0] r2_ror32_11_171_1094;
  reg  [31:0] arg_202_1096;
  reg  [31:0] r1_ror32_25_203_1100;
  reg  [24:0] r3_ror32_25_204_1097;
  reg  [6:0] r6_ror32_25_205_1098;
  reg  [31:0] r2_ror32_25_206_1099;
  reg  [31:0] x_22_1079;
  reg  [31:0] r1_e1_23_1085;
  reg  [31:0] r4_e1_24_1080;
  reg  [31:0] r6_e1_25_1081;
  reg  [31:0] r3_e1_26_1082;
  reg  [31:0] r8_e1_27_1083;
  reg  [31:0] r2_e1_28_1084;
  reg  [31:0] x_0_1104;
  reg  [31:0] y_1_1101;
  reg  [31:0] z_2_1102;
  reg  [31:0] r3_Ch_3_1107;
  reg  [31:0] r6_Ch_4_1103;
  reg  [31:0] r5_Ch_5_1105;
  reg  [31:0] r4_Ch_6_1106;
  reg  [31:0] arg_192_1115;
  reg  [31:0] r1_ror32_2_193_1119;
  reg  [1:0] r3_ror32_2_194_1116;
  reg  [29:0] r6_ror32_2_195_1117;
  reg  [31:0] r2_ror32_2_196_1118;
  reg  [31:0] arg_172_1120;
  reg  [31:0] r1_ror32_13_173_1124;
  reg  [12:0] r3_ror32_13_174_1121;
  reg  [18:0] r6_ror32_13_175_1122;
  reg  [31:0] r2_ror32_13_176_1123;
  reg  [31:0] arg_197_1125;
  reg  [31:0] r1_ror32_22_198_1129;
  reg  [21:0] r3_ror32_22_199_1126;
  reg  [9:0] r6_ror32_22_200_1127;
  reg  [31:0] r2_ror32_22_201_1128;
  reg  [31:0] x_15_1108;
  reg  [31:0] r1_e0_16_1114;
  reg  [31:0] r4_e0_17_1109;
  reg  [31:0] r6_e0_18_1110;
  reg  [31:0] r3_e0_19_1111;
  reg  [31:0] r8_e0_20_1112;
  reg  [31:0] r2_e0_21_1113;
  reg  [31:0] x_7_1130;
  reg  [31:0] y_8_1131;
  reg  [31:0] z_9_1134;
  reg  [31:0] r3_Maj_10_1137;
  reg  [31:0] r5_Maj_11_1132;
  reg  [31:0] r7_Maj_12_1133;
  reg  [31:0] r6_Maj_13_1135;
  reg  [31:0] r4_Maj_14_1136;
  reg  [31:0] arg_207_1145;
  reg  [31:0] r1_ror32_6_208_1149;
  reg  [5:0] r3_ror32_6_209_1146;
  reg  [25:0] r6_ror32_6_210_1147;
  reg  [31:0] r2_ror32_6_211_1148;
  reg  [31:0] arg_167_1150;
  reg  [31:0] r1_ror32_11_168_1154;
  reg  [10:0] r3_ror32_11_169_1151;
  reg  [20:0] r6_ror32_11_170_1152;
  reg  [31:0] r2_ror32_11_171_1153;
  reg  [31:0] arg_202_1155;
  reg  [31:0] r1_ror32_25_203_1159;
  reg  [24:0] r3_ror32_25_204_1156;
  reg  [6:0] r6_ror32_25_205_1157;
  reg  [31:0] r2_ror32_25_206_1158;
  reg  [31:0] x_22_1138;
  reg  [31:0] r1_e1_23_1144;
  reg  [31:0] r4_e1_24_1139;
  reg  [31:0] r6_e1_25_1140;
  reg  [31:0] r3_e1_26_1141;
  reg  [31:0] r8_e1_27_1142;
  reg  [31:0] r2_e1_28_1143;
  reg  [31:0] x_0_1163;
  reg  [31:0] y_1_1160;
  reg  [31:0] z_2_1161;
  reg  [31:0] r3_Ch_3_1166;
  reg  [31:0] r6_Ch_4_1162;
  reg  [31:0] r5_Ch_5_1164;
  reg  [31:0] r4_Ch_6_1165;
  reg  [31:0] arg_192_1174;
  reg  [31:0] r1_ror32_2_193_1178;
  reg  [1:0] r3_ror32_2_194_1175;
  reg  [29:0] r6_ror32_2_195_1176;
  reg  [31:0] r2_ror32_2_196_1177;
  reg  [31:0] arg_172_1179;
  reg  [31:0] r1_ror32_13_173_1183;
  reg  [12:0] r3_ror32_13_174_1180;
  reg  [18:0] r6_ror32_13_175_1181;
  reg  [31:0] r2_ror32_13_176_1182;
  reg  [31:0] arg_197_1184;
  reg  [31:0] r1_ror32_22_198_1188;
  reg  [21:0] r3_ror32_22_199_1185;
  reg  [9:0] r6_ror32_22_200_1186;
  reg  [31:0] r2_ror32_22_201_1187;
  reg  [31:0] x_15_1167;
  reg  [31:0] r1_e0_16_1173;
  reg  [31:0] r4_e0_17_1168;
  reg  [31:0] r6_e0_18_1169;
  reg  [31:0] r3_e0_19_1170;
  reg  [31:0] r8_e0_20_1171;
  reg  [31:0] r2_e0_21_1172;
  reg  [31:0] x_7_1189;
  reg  [31:0] y_8_1190;
  reg  [31:0] z_9_1193;
  reg  [31:0] r3_Maj_10_1196;
  reg  [31:0] r5_Maj_11_1191;
  reg  [31:0] r7_Maj_12_1192;
  reg  [31:0] r6_Maj_13_1194;
  reg  [31:0] r4_Maj_14_1195;
  reg  [31:0] a_30_602;
  reg  [31:0] b_31_604;
  reg  [31:0] c_32_605;
  reg  [31:0] r39_iterate_61_611;
  reg  [31:0] r188_iterate_150_700;
  reg  [31:0] d_33_609;
  reg  [31:0] e_34_588;
  reg  [31:0] f_35_592;
  reg  [31:0] g_36_593;
  reg  [31:0] h_37_590;
  reg  [31:0] idx_38_596;
  reg  [31:0] r9_iterate_39_717;
  reg  [31:0] r10_iterate_40_718;
  reg  [31:0] r11_iterate_41_719;
  reg  [31:0] r12_iterate_42_720;
  reg  [31:0] r13_iterate_43_721;
  reg  [31:0] r14_iterate_44_722;
  reg  [31:0] r15_iterate_45_723;
  reg  [31:0] r16_iterate_46_724;
  reg  [31:0] r23_iterate_47_589;
  reg  [31:0] r22_iterate_48_591;
  reg  [31:0] r25_iterate_49_594;
  reg  [31:0] r21_iterate_50_595;
  reg  [31:0] r27_iterate_51_597;
  reg  [31:0] r20_iterate_52_598;
  reg  [31:0] r30_iterate_53_599;
  reg  [31:0] r19_iterate_54_600;
  reg  [31:0] r17_iterate_55_601;
  reg  [31:0] r34_iterate_56_603;
  reg  [31:0] r36_iterate_57_606;
  reg  [31:0] r33_iterate_58_607;
  reg  [31:0] r18_iterate_59_608;
  reg  [31:0] r38_iterate_60_610;
  reg  [31:0] r133_iterate_119_669;
  reg  [31:0] r44_iterate_62_612;
  reg  [31:0] r69_iterate_77_627;
  reg  [31:0] r43_iterate_63_613;
  reg  [31:0] r46_iterate_64_614;
  reg  [31:0] r42_iterate_65_615;
  reg  [31:0] r48_iterate_66_616;
  reg  [31:0] r50_iterate_67_617;
  reg  [31:0] r41_iterate_68_618;
  reg  [31:0] r53_iterate_69_619;
  reg  [31:0] r55_iterate_70_620;
  reg  [31:0] r40_iterate_71_621;
  reg  [31:0] r59_iterate_72_622;
  reg  [31:0] r61_iterate_73_623;
  reg  [31:0] r148_iterate_126_676;
  reg  [31:0] r58_iterate_74_624;
  reg  [31:0] r63_iterate_75_625;
  reg  [31:0] r64_iterate_76_626;
  reg  [31:0] r119_iterate_107_657;
  reg  [31:0] r68_iterate_78_628;
  reg  [31:0] r71_iterate_79_629;
  reg  [31:0] r67_iterate_80_630;
  reg  [31:0] r73_iterate_81_631;
  reg  [31:0] r75_iterate_82_632;
  reg  [31:0] r66_iterate_83_633;
  reg  [31:0] r78_iterate_84_634;
  reg  [31:0] r80_iterate_85_635;
  reg  [31:0] r65_iterate_86_636;
  reg  [31:0] r84_iterate_87_637;
  reg  [31:0] r86_iterate_88_638;
  reg  [31:0] r83_iterate_89_639;
  reg  [31:0] r88_iterate_90_640;
  reg  [31:0] r89_iterate_91_641;
  reg  [31:0] r94_iterate_92_642;
  reg  [31:0] r93_iterate_93_643;
  reg  [31:0] r96_iterate_94_644;
  reg  [31:0] r92_iterate_95_645;
  reg  [31:0] r98_iterate_96_646;
  reg  [31:0] r100_iterate_97_647;
  reg  [31:0] r91_iterate_98_648;
  reg  [31:0] r103_iterate_99_649;
  reg  [31:0] r105_iterate_100_650;
  reg  [31:0] r90_iterate_101_651;
  reg  [31:0] r109_iterate_102_652;
  reg  [31:0] r111_iterate_103_653;
  reg  [31:0] r108_iterate_104_654;
  reg  [31:0] r113_iterate_105_655;
  reg  [31:0] r114_iterate_106_656;
  reg  [31:0] r213_iterate_165_715;
  reg  [31:0] r118_iterate_108_658;
  reg  [31:0] r121_iterate_109_659;
  reg  [31:0] r117_iterate_110_660;
  reg  [31:0] r123_iterate_111_661;
  reg  [31:0] r125_iterate_112_662;
  reg  [31:0] r116_iterate_113_663;
  reg  [31:0] r128_iterate_114_664;
  reg  [31:0] r130_iterate_115_665;
  reg  [31:0] r115_iterate_116_666;
  reg  [31:0] r134_iterate_117_667;
  reg  [31:0] r136_iterate_118_668;
  reg  [31:0] r138_iterate_120_670;
  reg  [31:0] r139_iterate_121_671;
  reg  [31:0] r144_iterate_122_672;
  reg  [31:0] r143_iterate_123_673;
  reg  [31:0] r146_iterate_124_674;
  reg  [31:0] r142_iterate_125_675;
  reg  [31:0] r150_iterate_127_677;
  reg  [31:0] r141_iterate_128_678;
  reg  [31:0] r153_iterate_129_679;
  reg  [31:0] r155_iterate_130_680;
  reg  [31:0] r140_iterate_131_681;
  reg  [31:0] r159_iterate_132_682;
  reg  [31:0] r161_iterate_133_683;
  reg  [31:0] r158_iterate_134_684;
  reg  [31:0] r163_iterate_135_685;
  reg  [31:0] r164_iterate_136_686;
  reg  [31:0] r169_iterate_137_687;
  reg  [31:0] r168_iterate_138_688;
  reg  [31:0] r171_iterate_139_689;
  reg  [31:0] r167_iterate_140_690;
  reg  [31:0] r173_iterate_141_691;
  reg  [31:0] r175_iterate_142_692;
  reg  [31:0] r166_iterate_143_693;
  reg  [31:0] r178_iterate_144_694;
  reg  [31:0] r180_iterate_145_695;
  reg  [31:0] r165_iterate_146_696;
  reg  [31:0] r184_iterate_147_697;
  reg  [31:0] r186_iterate_148_698;
  reg  [31:0] r183_iterate_149_699;
  reg  [31:0] r189_iterate_151_701;
  reg  [31:0] r194_iterate_152_702;
  reg  [31:0] r193_iterate_153_703;
  reg  [31:0] r196_iterate_154_704;
  reg  [31:0] r192_iterate_155_705;
  reg  [31:0] r198_iterate_156_706;
  reg  [31:0] r200_iterate_157_707;
  reg  [31:0] r191_iterate_158_708;
  reg  [31:0] r203_iterate_159_709;
  reg  [31:0] r205_iterate_160_710;
  reg  [31:0] r190_iterate_161_711;
  reg  [31:0] r209_iterate_162_712;
  reg  [31:0] r211_iterate_163_713;
  reg  [31:0] r208_iterate_164_714;
  reg  [31:0] r214_iterate_166_716;
  reg  [31:0] r__332_553;
  reg  [31:0] r0_transform_333_494;
  reg  r3_transform_334_495;
  reg  [31:0] r5_transform_335_496;
  reg  [31:0] r1_transform_336_497;
  reg  [7:0] r11_transform_337_498;
  reg  [7:0] r14_transform_338_499;
  reg  [15:0] r10_transform_339_500;
  reg  [7:0] r17_transform_340_501;
  reg  [23:0] r9_transform_341_502;
  reg  [7:0] r20_transform_342_503;
  reg  [31:0] r8_transform_343_504;
  reg  r26_transform_344_505;
  reg  [31:0] r33_transform_345_506;
  reg  [31:0] r35_transform_346_507;
  reg  [31:0] r31_transform_347_508;
  reg  [31:0] r38_transform_348_509;
  reg  [31:0] r40_transform_349_510;
  reg  [31:0] r30_transform_350_511;
  reg  [31:0] r45_transform_351_512;
  reg  [31:0] r47_transform_352_513;
  reg  [31:0] r43_transform_353_514;
  reg  [31:0] r29_transform_354_515;
  reg  [31:0] r50_transform_355_516;
  reg  [31:0] r52_transform_356_517;
  reg  [31:0] r28_transform_357_518;
  reg  [31:0] r66_transform_358_519;
  reg  [31:0] r57_transform_359_520;
  reg  [31:0] r70_transform_360_521;
  reg  [31:0] r58_transform_361_522;
  reg  [31:0] r74_transform_362_523;
  reg  [31:0] r59_transform_363_524;
  reg  [31:0] r78_transform_364_525;
  reg  [31:0] r60_transform_365_526;
  reg  [31:0] r82_transform_366_527;
  reg  [31:0] r61_transform_367_528;
  reg  [31:0] r86_transform_368_529;
  reg  [31:0] r62_transform_369_530;
  reg  [31:0] r90_transform_370_531;
  reg  [31:0] r63_transform_371_532;
  reg  [31:0] r94_transform_372_533;
  reg  [31:0] r64_transform_373_534;
  reg  r98_transform_374_535;
  reg  [31:0] r102_transform_375_536;
  reg  [31:0] r104_transform_376_537;
  reg  [31:0] r107_transform_377_538;
  reg  [31:0] r112_transform_378_539;
  reg  [31:0] r115_transform_379_540;
  reg  [31:0] r120_transform_380_541;
  reg  [31:0] r123_transform_381_542;
  reg  [31:0] r128_transform_382_543;
  reg  [31:0] r131_transform_383_544;
  reg  [31:0] r136_transform_384_545;
  reg  [31:0] r139_transform_385_546;
  reg  [31:0] r144_transform_386_547;
  reg  [31:0] r147_transform_387_548;
  reg  [31:0] r152_transform_388_549;
  reg  [31:0] r155_transform_389_550;
  reg  [31:0] r160_transform_390_551;
  reg  [31:0] r163_transform_391_552;
  reg  [15:0] r47_sha256_241_401;
  reg  [159:0] r29_sha256_295_455;
  reg  [31:0] r190_sha256_296_456;
  reg  [31:0] addr_231_392;
  reg  [31:0] blocks_232_393;
  reg  [255:0] r2_sha256_233_492;
  reg  [31:0] r5_sha256_234_394;
  reg  r7_sha256_235_395;
  reg  [31:0] r16_sha256_236_396;
  reg  [31:0] r50_sha256_237_397;
  reg  [7:0] r48_sha256_238_398;
  reg  [31:0] r57_sha256_239_399;
  reg  [7:0] r55_sha256_240_400;
  reg  [7:0] r237_sha256_318_478;
  reg  [31:0] r64_sha256_242_402;
  reg  [7:0] r62_sha256_243_403;
  reg  [23:0] r46_sha256_244_404;
  reg  [31:0] r71_sha256_245_405;
  reg  [7:0] r69_sha256_246_406;
  reg  [31:0] r45_sha256_247_407;
  reg  [31:0] r78_sha256_248_408;
  reg  [7:0] r76_sha256_249_409;
  reg  [39:0] r44_sha256_250_410;
  reg  [31:0] r85_sha256_251_411;
  reg  [7:0] r83_sha256_252_412;
  reg  [47:0] r43_sha256_253_413;
  reg  [31:0] r92_sha256_254_414;
  reg  [7:0] r90_sha256_255_415;
  reg  [55:0] r42_sha256_256_416;
  reg  [31:0] r99_sha256_257_417;
  reg  [7:0] r97_sha256_258_418;
  reg  [63:0] r41_sha256_259_419;
  reg  [31:0] r106_sha256_260_420;
  reg  [7:0] r104_sha256_261_421;
  reg  [71:0] r40_sha256_262_422;
  reg  [31:0] r113_sha256_263_423;
  reg  [7:0] r111_sha256_264_424;
  reg  [79:0] r39_sha256_265_425;
  reg  [31:0] r120_sha256_266_426;
  reg  [7:0] r118_sha256_267_427;
  reg  [87:0] r38_sha256_268_428;
  reg  [31:0] r127_sha256_269_429;
  reg  [7:0] r125_sha256_270_430;
  reg  [95:0] r37_sha256_271_431;
  reg  [31:0] r134_sha256_272_432;
  reg  [7:0] r132_sha256_273_433;
  reg  [103:0] r36_sha256_274_434;
  reg  [31:0] r141_sha256_275_435;
  reg  [7:0] r251_sha256_324_484;
  reg  [7:0] r139_sha256_276_436;
  reg  [111:0] r35_sha256_277_437;
  reg  [31:0] r148_sha256_278_438;
  reg  [7:0] r146_sha256_279_439;
  reg  [119:0] r34_sha256_280_440;
  reg  [31:0] r155_sha256_281_441;
  reg  [7:0] r153_sha256_282_442;
  reg  [127:0] r33_sha256_283_443;
  reg  [31:0] r162_sha256_284_444;
  reg  [7:0] r160_sha256_285_445;
  reg  [135:0] r32_sha256_286_446;
  reg  [31:0] r169_sha256_287_447;
  reg  [7:0] r167_sha256_288_448;
  reg  [143:0] r31_sha256_289_449;
  reg  [31:0] r176_sha256_290_450;
  reg  [7:0] r174_sha256_291_451;
  reg  [151:0] r30_sha256_292_452;
  reg  [31:0] r183_sha256_293_453;
  reg  [7:0] r181_sha256_294_454;
  reg  [7:0] r188_sha256_297_457;
  reg  [167:0] r28_sha256_298_458;
  reg  [31:0] r197_sha256_299_459;
  reg  [7:0] r195_sha256_300_460;
  reg  [175:0] r27_sha256_301_461;
  reg  [31:0] r204_sha256_302_462;
  reg  [7:0] r202_sha256_303_463;
  reg  [183:0] r26_sha256_304_464;
  reg  [31:0] r211_sha256_305_465;
  reg  [7:0] r209_sha256_306_466;
  reg  [191:0] r25_sha256_307_467;
  reg  [31:0] r218_sha256_308_468;
  reg  [7:0] r216_sha256_309_469;
  reg  [199:0] r24_sha256_310_470;
  reg  [31:0] r225_sha256_311_471;
  reg  [7:0] r223_sha256_312_472;
  reg  [207:0] r23_sha256_313_473;
  reg  [31:0] r232_sha256_314_474;
  reg  [7:0] r230_sha256_315_475;
  reg  [215:0] r22_sha256_316_476;
  reg  [31:0] r239_sha256_317_477;
  reg  [223:0] r21_sha256_319_479;
  reg  [31:0] r246_sha256_320_480;
  reg  [7:0] r244_sha256_321_481;
  reg  [231:0] r20_sha256_322_482;
  reg  [31:0] r253_sha256_323_483;
  reg  [239:0] r19_sha256_325_485;
  reg  [31:0] r260_sha256_326_486;
  reg  [7:0] r258_sha256_327_487;
  reg  [247:0] r18_sha256_328_488;
  reg  [31:0] r267_sha256_329_489;
  reg  [7:0] r265_sha256_330_490;
  reg  [255:0] r17_sha256_331_491;
  reg [31:0]  ext_task_arg_2_0;
  reg [31:0]  ext_task_arg_2_1;
  // Resources
  // add:16
  wire [31:0] add_16_s0;
  assign add_16_s0 = h_37_590;
  wire [31:0] add_16_s1;
  assign add_16_s1 = r23_iterate_47_589;
  wire [31:0] add_16_d0;
  assign add_16_d0 = add_16_s0 + add_16_s1;
  // add:17
  wire [31:0] add_17_s0;
  assign add_17_s0 = r22_iterate_48_591;
  wire [31:0] add_17_s1;
  assign add_17_s1 = r25_iterate_49_594;
  wire [31:0] add_17_d0;
  assign add_17_d0 = add_17_s0 + add_17_s1;
  // add:19
  wire [31:0] add_19_s0;
  assign add_19_s0 = r21_iterate_50_595;
  wire [31:0] add_19_s1;
  assign add_19_s1 = r27_iterate_51_597;
  wire [31:0] add_19_d0;
  assign add_19_d0 = add_19_s0 + add_19_s1;
  // add:21
  wire [31:0] add_21_s0;
  assign add_21_s0 = r20_iterate_52_598;
  wire [31:0] add_21_s1;
  assign add_21_s1 = r30_iterate_53_599;
  wire [31:0] add_21_d0;
  assign add_21_d0 = add_21_s0 + add_21_s1;
  // add:22
  wire [31:0] add_22_s0;
  assign add_22_s0 = r34_iterate_56_603;
  wire [31:0] add_22_s1;
  assign add_22_s1 = r36_iterate_57_606;
  wire [31:0] add_22_d0;
  assign add_22_d0 = add_22_s0 + add_22_s1;
  // add:23
  wire [31:0] add_23_s0;
  assign add_23_s0 = d_33_609;
  wire [31:0] add_23_s1;
  assign add_23_s1 = r17_iterate_55_601;
  wire [31:0] add_23_d0;
  assign add_23_d0 = add_23_s0 + add_23_s1;
  // add:24
  wire [31:0] add_24_s0;
  assign add_24_s0 = r17_iterate_55_601;
  wire [31:0] add_24_s1;
  assign add_24_s1 = r18_iterate_59_608;
  wire [31:0] add_24_d0;
  assign add_24_d0 = add_24_s0 + add_24_s1;
  // add:25
  wire [31:0] add_25_s0;
  assign add_25_s0 = g_36_593;
  wire [31:0] add_25_s1;
  assign add_25_s1 = r44_iterate_62_612;
  wire [31:0] add_25_d0;
  assign add_25_d0 = add_25_s0 + add_25_s1;
  // add:26
  wire [31:0] add_26_s0;
  assign add_26_s0 = r43_iterate_63_613;
  wire [31:0] add_26_s1;
  assign add_26_s1 = r46_iterate_64_614;
  wire [31:0] add_26_d0;
  assign add_26_d0 = add_26_s0 + add_26_s1;
  // add:27
  wire [31:0] add_27_s0;
  assign add_27_s0 = idx_38_596;
  wire [31:0] add_27_s1;
  assign add_27_s1 = 32'd1;
  wire [31:0] add_27_d0;
  assign add_27_d0 = add_27_s0 + add_27_s1;
  // add:28
  wire [31:0] add_28_s0;
  assign add_28_s0 = r42_iterate_65_615;
  wire [31:0] add_28_s1;
  assign add_28_s1 = r50_iterate_67_617;
  wire [31:0] add_28_d0;
  assign add_28_d0 = add_28_s0 + add_28_s1;
  // add:29
  wire [31:0] add_29_s0;
  assign add_29_s0 = idx_38_596;
  wire [31:0] add_29_s1;
  assign add_29_s1 = 32'd1;
  wire [31:0] add_29_d0;
  assign add_29_d0 = add_29_s0 + add_29_s1;
  // add:30
  wire [31:0] add_30_s0;
  assign add_30_s0 = r41_iterate_68_618;
  wire [31:0] add_30_s1;
  assign add_30_s1 = r55_iterate_70_620;
  wire [31:0] add_30_d0;
  assign add_30_d0 = add_30_s0 + add_30_s1;
  // add:31
  wire [31:0] add_31_s0;
  assign add_31_s0 = r59_iterate_72_622;
  wire [31:0] add_31_s1;
  assign add_31_s1 = r61_iterate_73_623;
  wire [31:0] add_31_d0;
  assign add_31_d0 = add_31_s0 + add_31_s1;
  // add:32
  wire [31:0] add_32_s0;
  assign add_32_s0 = c_32_605;
  wire [31:0] add_32_s1;
  assign add_32_s1 = r17_iterate_55_601;
  wire [31:0] add_32_d0;
  assign add_32_d0 = add_32_s0 + add_32_s1;
  // add:33
  wire [31:0] add_33_s0;
  assign add_33_s0 = r17_iterate_55_601;
  wire [31:0] add_33_s1;
  assign add_33_s1 = r18_iterate_59_608;
  wire [31:0] add_33_d0;
  assign add_33_d0 = add_33_s0 + add_33_s1;
  // add:34
  wire [31:0] add_34_s0;
  assign add_34_s0 = f_35_592;
  wire [31:0] add_34_s1;
  assign add_34_s1 = r69_iterate_77_627;
  wire [31:0] add_34_d0;
  assign add_34_d0 = add_34_s0 + add_34_s1;
  // add:35
  wire [31:0] add_35_s0;
  assign add_35_s0 = r68_iterate_78_628;
  wire [31:0] add_35_s1;
  assign add_35_s1 = r71_iterate_79_629;
  wire [31:0] add_35_d0;
  assign add_35_d0 = add_35_s0 + add_35_s1;
  // add:36
  wire [31:0] add_36_s0;
  assign add_36_s0 = idx_38_596;
  wire [31:0] add_36_s1;
  assign add_36_s1 = 32'd2;
  wire [31:0] add_36_d0;
  assign add_36_d0 = add_36_s0 + add_36_s1;
  // add:37
  wire [31:0] add_37_s0;
  assign add_37_s0 = r67_iterate_80_630;
  wire [31:0] add_37_s1;
  assign add_37_s1 = r75_iterate_82_632;
  wire [31:0] add_37_d0;
  assign add_37_d0 = add_37_s0 + add_37_s1;
  // add:38
  wire [31:0] add_38_s0;
  assign add_38_s0 = idx_38_596;
  wire [31:0] add_38_s1;
  assign add_38_s1 = 32'd2;
  wire [31:0] add_38_d0;
  assign add_38_d0 = add_38_s0 + add_38_s1;
  // add:39
  wire [31:0] add_39_s0;
  assign add_39_s0 = r66_iterate_83_633;
  wire [31:0] add_39_s1;
  assign add_39_s1 = r80_iterate_85_635;
  wire [31:0] add_39_d0;
  assign add_39_d0 = add_39_s0 + add_39_s1;
  // add:40
  wire [31:0] add_40_s0;
  assign add_40_s0 = r84_iterate_87_637;
  wire [31:0] add_40_s1;
  assign add_40_s1 = r86_iterate_88_638;
  wire [31:0] add_40_d0;
  assign add_40_d0 = add_40_s0 + add_40_s1;
  // add:41
  wire [31:0] add_41_s0;
  assign add_41_s0 = b_31_604;
  wire [31:0] add_41_s1;
  assign add_41_s1 = r17_iterate_55_601;
  wire [31:0] add_41_d0;
  assign add_41_d0 = add_41_s0 + add_41_s1;
  // add:42
  wire [31:0] add_42_s0;
  assign add_42_s0 = r17_iterate_55_601;
  wire [31:0] add_42_s1;
  assign add_42_s1 = r18_iterate_59_608;
  wire [31:0] add_42_d0;
  assign add_42_d0 = add_42_s0 + add_42_s1;
  // add:43
  wire [31:0] add_43_s0;
  assign add_43_s0 = e_34_588;
  wire [31:0] add_43_s1;
  assign add_43_s1 = r94_iterate_92_642;
  wire [31:0] add_43_d0;
  assign add_43_d0 = add_43_s0 + add_43_s1;
  // add:44
  wire [31:0] add_44_s0;
  assign add_44_s0 = r93_iterate_93_643;
  wire [31:0] add_44_s1;
  assign add_44_s1 = r96_iterate_94_644;
  wire [31:0] add_44_d0;
  assign add_44_d0 = add_44_s0 + add_44_s1;
  // add:45
  wire [31:0] add_45_s0;
  assign add_45_s0 = idx_38_596;
  wire [31:0] add_45_s1;
  assign add_45_s1 = 32'd3;
  wire [31:0] add_45_d0;
  assign add_45_d0 = add_45_s0 + add_45_s1;
  // add:46
  wire [31:0] add_46_s0;
  assign add_46_s0 = r92_iterate_95_645;
  wire [31:0] add_46_s1;
  assign add_46_s1 = r100_iterate_97_647;
  wire [31:0] add_46_d0;
  assign add_46_d0 = add_46_s0 + add_46_s1;
  // add:47
  wire [31:0] add_47_s0;
  assign add_47_s0 = idx_38_596;
  wire [31:0] add_47_s1;
  assign add_47_s1 = 32'd3;
  wire [31:0] add_47_d0;
  assign add_47_d0 = add_47_s0 + add_47_s1;
  // add:48
  wire [31:0] add_48_s0;
  assign add_48_s0 = r91_iterate_98_648;
  wire [31:0] add_48_s1;
  assign add_48_s1 = r105_iterate_100_650;
  wire [31:0] add_48_d0;
  assign add_48_d0 = add_48_s0 + add_48_s1;
  // add:49
  wire [31:0] add_49_s0;
  assign add_49_s0 = r109_iterate_102_652;
  wire [31:0] add_49_s1;
  assign add_49_s1 = r111_iterate_103_653;
  wire [31:0] add_49_d0;
  assign add_49_d0 = add_49_s0 + add_49_s1;
  // add:50
  wire [31:0] add_50_s0;
  assign add_50_s0 = a_30_602;
  wire [31:0] add_50_s1;
  assign add_50_s1 = r17_iterate_55_601;
  wire [31:0] add_50_d0;
  assign add_50_d0 = add_50_s0 + add_50_s1;
  // add:51
  wire [31:0] add_51_s0;
  assign add_51_s0 = r17_iterate_55_601;
  wire [31:0] add_51_s1;
  assign add_51_s1 = r18_iterate_59_608;
  wire [31:0] add_51_d0;
  assign add_51_d0 = add_51_s0 + add_51_s1;
  // add:52
  wire [31:0] add_52_s0;
  assign add_52_s0 = d_33_609;
  wire [31:0] add_52_s1;
  assign add_52_s1 = r119_iterate_107_657;
  wire [31:0] add_52_d0;
  assign add_52_d0 = add_52_s0 + add_52_s1;
  // add:53
  wire [31:0] add_53_s0;
  assign add_53_s0 = r118_iterate_108_658;
  wire [31:0] add_53_s1;
  assign add_53_s1 = r121_iterate_109_659;
  wire [31:0] add_53_d0;
  assign add_53_d0 = add_53_s0 + add_53_s1;
  // add:54
  wire [31:0] add_54_s0;
  assign add_54_s0 = idx_38_596;
  wire [31:0] add_54_s1;
  assign add_54_s1 = 32'd4;
  wire [31:0] add_54_d0;
  assign add_54_d0 = add_54_s0 + add_54_s1;
  // add:55
  wire [31:0] add_55_s0;
  assign add_55_s0 = r117_iterate_110_660;
  wire [31:0] add_55_s1;
  assign add_55_s1 = r125_iterate_112_662;
  wire [31:0] add_55_d0;
  assign add_55_d0 = add_55_s0 + add_55_s1;
  // add:56
  wire [31:0] add_56_s0;
  assign add_56_s0 = idx_38_596;
  wire [31:0] add_56_s1;
  assign add_56_s1 = 32'd4;
  wire [31:0] add_56_d0;
  assign add_56_d0 = add_56_s0 + add_56_s1;
  // add:57
  wire [31:0] add_57_s0;
  assign add_57_s0 = r116_iterate_113_663;
  wire [31:0] add_57_s1;
  assign add_57_s1 = r130_iterate_115_665;
  wire [31:0] add_57_d0;
  assign add_57_d0 = add_57_s0 + add_57_s1;
  // add:58
  wire [31:0] add_58_s0;
  assign add_58_s0 = r134_iterate_117_667;
  wire [31:0] add_58_s1;
  assign add_58_s1 = r136_iterate_118_668;
  wire [31:0] add_58_d0;
  assign add_58_d0 = add_58_s0 + add_58_s1;
  // add:59
  wire [31:0] add_59_s0;
  assign add_59_s0 = h_37_590;
  wire [31:0] add_59_s1;
  assign add_59_s1 = r17_iterate_55_601;
  wire [31:0] add_59_d0;
  assign add_59_d0 = add_59_s0 + add_59_s1;
  // add:60
  wire [31:0] add_60_s0;
  assign add_60_s0 = r17_iterate_55_601;
  wire [31:0] add_60_s1;
  assign add_60_s1 = r18_iterate_59_608;
  wire [31:0] add_60_d0;
  assign add_60_d0 = add_60_s0 + add_60_s1;
  // add:61
  wire [31:0] add_61_s0;
  assign add_61_s0 = c_32_605;
  wire [31:0] add_61_s1;
  assign add_61_s1 = r144_iterate_122_672;
  wire [31:0] add_61_d0;
  assign add_61_d0 = add_61_s0 + add_61_s1;
  // add:62
  wire [31:0] add_62_s0;
  assign add_62_s0 = r143_iterate_123_673;
  wire [31:0] add_62_s1;
  assign add_62_s1 = r146_iterate_124_674;
  wire [31:0] add_62_d0;
  assign add_62_d0 = add_62_s0 + add_62_s1;
  // add:63
  wire [31:0] add_63_s0;
  assign add_63_s0 = idx_38_596;
  wire [31:0] add_63_s1;
  assign add_63_s1 = 32'd5;
  wire [31:0] add_63_d0;
  assign add_63_d0 = add_63_s0 + add_63_s1;
  // add:64
  wire [31:0] add_64_s0;
  assign add_64_s0 = r142_iterate_125_675;
  wire [31:0] add_64_s1;
  assign add_64_s1 = r150_iterate_127_677;
  wire [31:0] add_64_d0;
  assign add_64_d0 = add_64_s0 + add_64_s1;
  // add:65
  wire [31:0] add_65_s0;
  assign add_65_s0 = idx_38_596;
  wire [31:0] add_65_s1;
  assign add_65_s1 = 32'd5;
  wire [31:0] add_65_d0;
  assign add_65_d0 = add_65_s0 + add_65_s1;
  // add:66
  wire [31:0] add_66_s0;
  assign add_66_s0 = r141_iterate_128_678;
  wire [31:0] add_66_s1;
  assign add_66_s1 = r155_iterate_130_680;
  wire [31:0] add_66_d0;
  assign add_66_d0 = add_66_s0 + add_66_s1;
  // add:67
  wire [31:0] add_67_s0;
  assign add_67_s0 = r159_iterate_132_682;
  wire [31:0] add_67_s1;
  assign add_67_s1 = r161_iterate_133_683;
  wire [31:0] add_67_d0;
  assign add_67_d0 = add_67_s0 + add_67_s1;
  // add:68
  wire [31:0] add_68_s0;
  assign add_68_s0 = g_36_593;
  wire [31:0] add_68_s1;
  assign add_68_s1 = r17_iterate_55_601;
  wire [31:0] add_68_d0;
  assign add_68_d0 = add_68_s0 + add_68_s1;
  // add:69
  wire [31:0] add_69_s0;
  assign add_69_s0 = r17_iterate_55_601;
  wire [31:0] add_69_s1;
  assign add_69_s1 = r18_iterate_59_608;
  wire [31:0] add_69_d0;
  assign add_69_d0 = add_69_s0 + add_69_s1;
  // add:70
  wire [31:0] add_70_s0;
  assign add_70_s0 = b_31_604;
  wire [31:0] add_70_s1;
  assign add_70_s1 = r169_iterate_137_687;
  wire [31:0] add_70_d0;
  assign add_70_d0 = add_70_s0 + add_70_s1;
  // add:71
  wire [31:0] add_71_s0;
  assign add_71_s0 = r168_iterate_138_688;
  wire [31:0] add_71_s1;
  assign add_71_s1 = r171_iterate_139_689;
  wire [31:0] add_71_d0;
  assign add_71_d0 = add_71_s0 + add_71_s1;
  // add:72
  wire [31:0] add_72_s0;
  assign add_72_s0 = idx_38_596;
  wire [31:0] add_72_s1;
  assign add_72_s1 = 32'd6;
  wire [31:0] add_72_d0;
  assign add_72_d0 = add_72_s0 + add_72_s1;
  // add:73
  wire [31:0] add_73_s0;
  assign add_73_s0 = r167_iterate_140_690;
  wire [31:0] add_73_s1;
  assign add_73_s1 = r175_iterate_142_692;
  wire [31:0] add_73_d0;
  assign add_73_d0 = add_73_s0 + add_73_s1;
  // add:74
  wire [31:0] add_74_s0;
  assign add_74_s0 = idx_38_596;
  wire [31:0] add_74_s1;
  assign add_74_s1 = 32'd6;
  wire [31:0] add_74_d0;
  assign add_74_d0 = add_74_s0 + add_74_s1;
  // add:75
  wire [31:0] add_75_s0;
  assign add_75_s0 = r166_iterate_143_693;
  wire [31:0] add_75_s1;
  assign add_75_s1 = r180_iterate_145_695;
  wire [31:0] add_75_d0;
  assign add_75_d0 = add_75_s0 + add_75_s1;
  // add:76
  wire [31:0] add_76_s0;
  assign add_76_s0 = r184_iterate_147_697;
  wire [31:0] add_76_s1;
  assign add_76_s1 = r186_iterate_148_698;
  wire [31:0] add_76_d0;
  assign add_76_d0 = add_76_s0 + add_76_s1;
  // add:77
  wire [31:0] add_77_s0;
  assign add_77_s0 = f_35_592;
  wire [31:0] add_77_s1;
  assign add_77_s1 = r17_iterate_55_601;
  wire [31:0] add_77_d0;
  assign add_77_d0 = add_77_s0 + add_77_s1;
  // add:78
  wire [31:0] add_78_s0;
  assign add_78_s0 = r17_iterate_55_601;
  wire [31:0] add_78_s1;
  assign add_78_s1 = r18_iterate_59_608;
  wire [31:0] add_78_d0;
  assign add_78_d0 = add_78_s0 + add_78_s1;
  // add:79
  wire [31:0] add_79_s0;
  assign add_79_s0 = a_30_602;
  wire [31:0] add_79_s1;
  assign add_79_s1 = r194_iterate_152_702;
  wire [31:0] add_79_d0;
  assign add_79_d0 = add_79_s0 + add_79_s1;
  // add:80
  wire [31:0] add_80_s0;
  assign add_80_s0 = r193_iterate_153_703;
  wire [31:0] add_80_s1;
  assign add_80_s1 = r196_iterate_154_704;
  wire [31:0] add_80_d0;
  assign add_80_d0 = add_80_s0 + add_80_s1;
  // add:81
  wire [31:0] add_81_s0;
  assign add_81_s0 = idx_38_596;
  wire [31:0] add_81_s1;
  assign add_81_s1 = 32'd7;
  wire [31:0] add_81_d0;
  assign add_81_d0 = add_81_s0 + add_81_s1;
  // add:82
  wire [31:0] add_82_s0;
  assign add_82_s0 = r192_iterate_155_705;
  wire [31:0] add_82_s1;
  assign add_82_s1 = r200_iterate_157_707;
  wire [31:0] add_82_d0;
  assign add_82_d0 = add_82_s0 + add_82_s1;
  // add:83
  wire [31:0] add_83_s0;
  assign add_83_s0 = idx_38_596;
  wire [31:0] add_83_s1;
  assign add_83_s1 = 32'd7;
  wire [31:0] add_83_d0;
  assign add_83_d0 = add_83_s0 + add_83_s1;
  // add:84
  wire [31:0] add_84_s0;
  assign add_84_s0 = r191_iterate_158_708;
  wire [31:0] add_84_s1;
  assign add_84_s1 = r205_iterate_160_710;
  wire [31:0] add_84_d0;
  assign add_84_d0 = add_84_s0 + add_84_s1;
  // add:85
  wire [31:0] add_85_s0;
  assign add_85_s0 = r209_iterate_162_712;
  wire [31:0] add_85_s1;
  assign add_85_s1 = r211_iterate_163_713;
  wire [31:0] add_85_d0;
  assign add_85_d0 = add_85_s0 + add_85_s1;
  // add:86
  wire [31:0] add_86_s0;
  assign add_86_s0 = e_34_588;
  wire [31:0] add_86_s1;
  assign add_86_s1 = r17_iterate_55_601;
  wire [31:0] add_86_d0;
  assign add_86_d0 = add_86_s0 + add_86_s1;
  // add:87
  wire [31:0] add_87_s0;
  assign add_87_s0 = r17_iterate_55_601;
  wire [31:0] add_87_s1;
  assign add_87_s1 = r18_iterate_59_608;
  wire [31:0] add_87_d0;
  assign add_87_d0 = add_87_s0 + add_87_s1;
  // gt:124
  wire [31:0] gt_124_s0;
  assign gt_124_s0 = blocks_232_393;
  wire [31:0] gt_124_s1;
  assign gt_124_s1 = r5_sha256_234_394;
  wire gt_124_d0;
  assign gt_124_d0 = gt_124_s0 > gt_124_s1;
  wire [3:0]  mem_1_2_125_p0_addr;
  wire [31:0]  mem_1_2_125_p0_rdata;
  wire [31:0]  mem_1_2_125_p0_wdata;
  wire mem_1_2_125_p0_wen;
  wire [3:0]  mem_1_2_125_p1_addr;
  wire [31:0]  mem_1_2_125_p1_rdata;
  wire [31:0]  mem_1_2_125_p1_wdata;
  wire mem_1_2_125_p1_wen;
  reg mem_1_2_125_1_2_125_ack;
  assign mem_1_2_125_p0_addr = mem_1_2_125_1_2_125_p0_addr;
  assign mem_1_2_125_p0_wdata = mem_1_2_125_1_2_125_p0_wdata;
  assign mem_1_2_125_p0_wen = (mem_1_2_125_1_2_125_p0_wen & !mem_1_2_125_1_2_125_ack);
  reg [3:0] mem_1_2_125_1_2_125_p0_addr;
  reg mem_1_2_125_1_2_125_req;
  reg [31:0] mem_1_2_125_1_2_125_p0_wdata;
  reg mem_1_2_125_1_2_125_p0_wen;
  reg [31:0] mem_1_2_125_1_2_125_rbuf;
  reg [31:0] axi_addr2_126;
  reg axi_wen2_126;
  reg axi_req2_126;
  wire axi_ack2_126;
  reg [3:0] axi_len2_126;
  reg [3:0] axi_start2_126;
  // add:127
  wire [31:0] add_127_s0;
  assign add_127_s0 = addr_231_392;
  wire [31:0] add_127_s1;
  assign add_127_s1 = 32'd64;
  wire [31:0] add_127_d0;
  assign add_127_d0 = add_127_s0 + add_127_s1;
  // add:128
  wire [31:0] add_128_s0;
  assign add_128_s0 = r5_sha256_234_394;
  wire [31:0] add_128_s1;
  assign add_128_s1 = 32'd1;
  wire [31:0] add_128_d0;
  assign add_128_d0 = add_128_s0 + add_128_s1;
  // gt:194
  wire [31:0] gt_194_s0;
  assign gt_194_s0 = 32'd16;
  wire [31:0] gt_194_s1;
  assign gt_194_s1 = r0_transform_333_494;
  wire gt_194_d0;
  assign gt_194_d0 = gt_194_s0 > gt_194_s1;
  // add:202
  wire [31:0] add_202_s0;
  assign add_202_s0 = r0_transform_333_494;
  wire [31:0] add_202_s1;
  assign add_202_s1 = 32'd1;
  wire [31:0] add_202_d0;
  assign add_202_d0 = add_202_s0 + add_202_s1;
  // gt:203
  wire [31:0] gt_203_s0;
  assign gt_203_s0 = 32'd64;
  wire [31:0] gt_203_s1;
  assign gt_203_s1 = r0_transform_333_494;
  wire gt_203_d0;
  assign gt_203_d0 = gt_203_s0 > gt_203_s1;
  // sub:204
  wire [31:0] sub_204_s0;
  assign sub_204_s0 = r0_transform_333_494;
  wire [31:0] sub_204_s1;
  assign sub_204_s1 = 32'd2;
  wire [31:0] sub_204_d0;
  assign sub_204_d0 = sub_204_s0 - sub_204_s1;
  // sub:205
  wire [31:0] sub_205_s0;
  assign sub_205_s0 = r0_transform_333_494;
  wire [31:0] sub_205_s1;
  assign sub_205_s1 = 32'd7;
  wire [31:0] sub_205_d0;
  assign sub_205_d0 = sub_205_s0 - sub_205_s1;
  // add:206
  wire [31:0] add_206_s0;
  assign add_206_s0 = r31_transform_347_508;
  wire [31:0] add_206_s1;
  assign add_206_s1 = r40_transform_349_510;
  wire [31:0] add_206_d0;
  assign add_206_d0 = add_206_s0 + add_206_s1;
  // sub:207
  wire [31:0] sub_207_s0;
  assign sub_207_s0 = r0_transform_333_494;
  wire [31:0] sub_207_s1;
  assign sub_207_s1 = 32'd15;
  wire [31:0] sub_207_d0;
  assign sub_207_d0 = sub_207_s0 - sub_207_s1;
  // add:208
  wire [31:0] add_208_s0;
  assign add_208_s0 = r30_transform_350_511;
  wire [31:0] add_208_s1;
  assign add_208_s1 = r43_transform_353_514;
  wire [31:0] add_208_d0;
  assign add_208_d0 = add_208_s0 + add_208_s1;
  // sub:209
  wire [31:0] sub_209_s0;
  assign sub_209_s0 = r0_transform_333_494;
  wire [31:0] sub_209_s1;
  assign sub_209_s1 = 32'd16;
  wire [31:0] sub_209_d0;
  assign sub_209_d0 = sub_209_s0 - sub_209_s1;
  // add:210
  wire [31:0] add_210_s0;
  assign add_210_s0 = r29_transform_354_515;
  wire [31:0] add_210_s1;
  assign add_210_s1 = r52_transform_356_517;
  wire [31:0] add_210_d0;
  assign add_210_d0 = add_210_s0 + add_210_s1;
  // add:211
  wire [31:0] add_211_s0;
  assign add_211_s0 = r0_transform_333_494;
  wire [31:0] add_211_s1;
  assign add_211_s1 = 32'd1;
  wire [31:0] add_211_d0;
  assign add_211_d0 = add_211_s0 + add_211_s1;
  // gt:212
  wire [31:0] gt_212_s0;
  assign gt_212_s0 = 32'd64;
  wire [31:0] gt_212_s1;
  assign gt_212_s1 = r0_transform_333_494;
  wire gt_212_d0;
  assign gt_212_d0 = gt_212_s0 > gt_212_s1;
  // add:213
  wire [31:0] add_213_s0;
  assign add_213_s0 = r0_transform_333_494;
  wire [31:0] add_213_s1;
  assign add_213_s1 = 32'd8;
  wire [31:0] add_213_d0;
  assign add_213_d0 = add_213_s0 + add_213_s1;
  // add:214
  wire [31:0] add_214_s0;
  assign add_214_s0 = r104_transform_376_537;
  wire [31:0] add_214_s1;
  assign add_214_s1 = r57_transform_359_520;
  wire [31:0] add_214_d0;
  assign add_214_d0 = add_214_s0 + add_214_s1;
  // add:215
  wire [31:0] add_215_s0;
  assign add_215_s0 = r112_transform_378_539;
  wire [31:0] add_215_s1;
  assign add_215_s1 = r58_transform_361_522;
  wire [31:0] add_215_d0;
  assign add_215_d0 = add_215_s0 + add_215_s1;
  // add:216
  wire [31:0] add_216_s0;
  assign add_216_s0 = r120_transform_380_541;
  wire [31:0] add_216_s1;
  assign add_216_s1 = r59_transform_363_524;
  wire [31:0] add_216_d0;
  assign add_216_d0 = add_216_s0 + add_216_s1;
  // add:217
  wire [31:0] add_217_s0;
  assign add_217_s0 = r128_transform_382_543;
  wire [31:0] add_217_s1;
  assign add_217_s1 = r60_transform_365_526;
  wire [31:0] add_217_d0;
  assign add_217_d0 = add_217_s0 + add_217_s1;
  // add:218
  wire [31:0] add_218_s0;
  assign add_218_s0 = r136_transform_384_545;
  wire [31:0] add_218_s1;
  assign add_218_s1 = r61_transform_367_528;
  wire [31:0] add_218_d0;
  assign add_218_d0 = add_218_s0 + add_218_s1;
  // add:219
  wire [31:0] add_219_s0;
  assign add_219_s0 = r144_transform_386_547;
  wire [31:0] add_219_s1;
  assign add_219_s1 = r62_transform_369_530;
  wire [31:0] add_219_d0;
  assign add_219_d0 = add_219_s0 + add_219_s1;
  // add:220
  wire [31:0] add_220_s0;
  assign add_220_s0 = r152_transform_388_549;
  wire [31:0] add_220_s1;
  assign add_220_s1 = r63_transform_371_532;
  wire [31:0] add_220_d0;
  assign add_220_d0 = add_220_s0 + add_220_s1;
  // add:221
  wire [31:0] add_221_s0;
  assign add_221_s0 = r160_transform_390_551;
  wire [31:0] add_221_s1;
  assign add_221_s1 = r64_transform_373_534;
  wire [31:0] add_221_d0;
  assign add_221_d0 = add_221_s0 + add_221_s1;
  reg [2:0] sram_addr_2;
  wire [31:0] sram_rdata_2;
  reg [31:0] sram_wdata_2;
  reg sram_wdata_en_2;
  reg [5:0] sram_addr_222;
  wire [31:0] sram_rdata_222;
  reg [31:0] sram_wdata_222;
  reg sram_wdata_en_222;
  reg [5:0] sram_addr_223;
  wire [31:0] sram_rdata_223;
  reg [31:0] sram_wdata_223;
  reg sram_wdata_en_223;
  // Insn wires
  wire  [31:0] insn_o_2_2_0;
  wire  [31:0] insn_o_2_2_1;
  wire  [31:0] insn_o_2_8_0;
  wire  insn_o_2_10_0;
  wire  [31:0] insn_o_2_25_0;
  wire  [31:0] insn_o_2_27_0;
  wire  [31:0] insn_o_2_29_0;
  wire  [31:0] insn_o_2_5_0;
  wire  [7:0] insn_o_2_39_0;
  wire  [31:0] insn_o_2_14_0;
  wire  [7:0] insn_o_2_48_0;
  wire  [15:0] insn_o_2_50_0;
  wire  [31:0] insn_o_2_19_0;
  wire  [7:0] insn_o_2_59_0;
  wire  [23:0] insn_o_2_61_0;
  wire  [31:0] insn_o_2_22_0;
  wire  [7:0] insn_o_2_70_0;
  wire  [31:0] insn_o_2_72_0;
  wire  [31:0] insn_o_2_31_0;
  wire  [7:0] insn_o_2_81_0;
  wire  [39:0] insn_o_2_83_0;
  wire  [31:0] insn_o_2_35_0;
  wire  [7:0] insn_o_2_92_0;
  wire  [47:0] insn_o_2_94_0;
  wire  [31:0] insn_o_2_41_0;
  wire  [7:0] insn_o_2_103_0;
  wire  [55:0] insn_o_2_105_0;
  wire  [31:0] insn_o_2_44_0;
  wire  [7:0] insn_o_2_114_0;
  wire  [63:0] insn_o_2_116_0;
  wire  [31:0] insn_o_2_52_0;
  wire  [7:0] insn_o_2_125_0;
  wire  [71:0] insn_o_2_127_0;
  wire  [31:0] insn_o_2_55_0;
  wire  [7:0] insn_o_2_136_0;
  wire  [79:0] insn_o_2_138_0;
  wire  [31:0] insn_o_2_63_0;
  wire  [7:0] insn_o_2_147_0;
  wire  [87:0] insn_o_2_149_0;
  wire  [31:0] insn_o_2_66_0;
  wire  [7:0] insn_o_2_158_0;
  wire  [95:0] insn_o_2_160_0;
  wire  [31:0] insn_o_2_74_0;
  wire  [7:0] insn_o_2_169_0;
  wire  [103:0] insn_o_2_171_0;
  wire  [31:0] insn_o_2_77_0;
  wire  [7:0] insn_o_2_180_0;
  wire  [111:0] insn_o_2_182_0;
  wire  [31:0] insn_o_2_85_0;
  wire  [7:0] insn_o_2_191_0;
  wire  [119:0] insn_o_2_193_0;
  wire  [31:0] insn_o_2_88_0;
  wire  [7:0] insn_o_2_202_0;
  wire  [127:0] insn_o_2_204_0;
  wire  [31:0] insn_o_2_96_0;
  wire  [7:0] insn_o_2_213_0;
  wire  [135:0] insn_o_2_215_0;
  wire  [31:0] insn_o_2_99_0;
  wire  [7:0] insn_o_2_224_0;
  wire  [143:0] insn_o_2_226_0;
  wire  [31:0] insn_o_2_107_0;
  wire  [7:0] insn_o_2_235_0;
  wire  [151:0] insn_o_2_237_0;
  wire  [31:0] insn_o_2_110_0;
  wire  [7:0] insn_o_2_246_0;
  wire  [159:0] insn_o_2_248_0;
  wire  [31:0] insn_o_2_118_0;
  wire  [7:0] insn_o_2_257_0;
  wire  [167:0] insn_o_2_259_0;
  wire  [31:0] insn_o_2_121_0;
  wire  [7:0] insn_o_2_268_0;
  wire  [175:0] insn_o_2_270_0;
  wire  [31:0] insn_o_2_129_0;
  wire  [7:0] insn_o_2_279_0;
  wire  [183:0] insn_o_2_281_0;
  wire  [31:0] insn_o_2_132_0;
  wire  [7:0] insn_o_2_290_0;
  wire  [191:0] insn_o_2_292_0;
  wire  [31:0] insn_o_2_140_0;
  wire  [7:0] insn_o_2_301_0;
  wire  [199:0] insn_o_2_303_0;
  wire  [31:0] insn_o_2_143_0;
  wire  [7:0] insn_o_2_312_0;
  wire  [207:0] insn_o_2_314_0;
  wire  [31:0] insn_o_2_151_0;
  wire  [7:0] insn_o_2_323_0;
  wire  [215:0] insn_o_2_325_0;
  wire  [31:0] insn_o_2_154_0;
  wire  [7:0] insn_o_2_334_0;
  wire  [223:0] insn_o_2_336_0;
  wire  [31:0] insn_o_2_162_0;
  wire  [7:0] insn_o_2_345_0;
  wire  [231:0] insn_o_2_347_0;
  wire  [31:0] insn_o_2_165_0;
  wire  [7:0] insn_o_2_356_0;
  wire  [239:0] insn_o_2_358_0;
  wire  [31:0] insn_o_2_173_0;
  wire  [7:0] insn_o_2_367_0;
  wire  [247:0] insn_o_2_369_0;
  wire  [31:0] insn_o_2_176_0;
  wire  [7:0] insn_o_2_378_0;
  wire  [255:0] insn_o_2_380_0;
  wire  [255:0] insn_o_2_382_0;
  wire  [31:0] insn_o_2_442_0;
  wire  insn_o_2_445_0;
  wire  [31:0] insn_o_2_450_0;
  wire  [31:0] insn_o_2_452_0;
  wire  [7:0] insn_o_2_456_0;
  wire  [7:0] insn_o_2_460_0;
  wire  [15:0] insn_o_2_462_0;
  wire  [7:0] insn_o_2_466_0;
  wire  [23:0] insn_o_2_468_0;
  wire  [7:0] insn_o_2_472_0;
  wire  [31:0] insn_o_2_474_0;
  wire  [31:0] insn_o_2_480_0;
  wire  [31:0] insn_o_2_484_0;
  wire  insn_o_2_487_0;
  wire  [31:0] insn_o_2_492_0;
  wire  [31:0] insn_o_2_198_0;
  wire  [31:0] insn_o_2_500_0;
  wire  [31:0] insn_o_2_502_0;
  wire  [31:0] insn_o_2_504_0;
  wire  [31:0] insn_o_2_206_0;
  wire  [31:0] insn_o_2_510_0;
  wire  [31:0] insn_o_2_514_0;
  wire  [31:0] insn_o_2_209_0;
  wire  [31:0] insn_o_2_522_0;
  wire  [31:0] insn_o_2_524_0;
  wire  [31:0] insn_o_2_525_0;
  wire  [31:0] insn_o_2_528_0;
  wire  [31:0] insn_o_2_217_0;
  wire  [31:0] insn_o_2_534_0;
  wire  [31:0] insn_o_2_540_0;
  wire  [31:0] insn_o_2_222_0;
  wire  [31:0] insn_o_2_548_0;
  wire  [31:0] insn_o_2_229_0;
  wire  [31:0] insn_o_2_555_0;
  wire  [31:0] insn_o_2_233_0;
  wire  [31:0] insn_o_2_562_0;
  wire  [31:0] insn_o_2_240_0;
  wire  [31:0] insn_o_2_569_0;
  wire  [31:0] insn_o_2_244_0;
  wire  [31:0] insn_o_2_576_0;
  wire  [31:0] insn_o_2_251_0;
  wire  [31:0] insn_o_2_583_0;
  wire  [31:0] insn_o_2_255_0;
  wire  [31:0] insn_o_2_590_0;
  wire  [31:0] insn_o_2_262_0;
  wire  [31:0] insn_o_2_597_0;
  wire  [31:0] insn_o_2_600_0;
  wire  insn_o_2_603_0;
  wire  [31:0] insn_o_2_609_0;
  wire  [31:0] insn_o_2_610_0;
  wire  [31:0] insn_o_2_611_0;
  wire  [31:0] insn_o_2_612_0;
  wire  [31:0] insn_o_2_613_0;
  wire  [31:0] insn_o_2_614_0;
  wire  [31:0] insn_o_2_615_0;
  wire  [31:0] insn_o_2_616_0;
  wire  [31:0] insn_o_2_617_0;
  wire  [31:0] insn_o_2_619_0;
  wire  [31:0] insn_o_2_620_0;
  wire  [31:0] insn_o_2_621_0;
  wire  [31:0] insn_o_2_622_0;
  wire  [31:0] insn_o_2_623_0;
  wire  [31:0] insn_o_2_624_0;
  wire  [31:0] insn_o_2_625_0;
  wire  [31:0] insn_o_2_626_0;
  wire  [31:0] insn_o_2_628_0;
  wire  [31:0] insn_o_2_630_0;
  wire  [31:0] insn_o_2_266_0;
  wire  [31:0] insn_o_2_638_0;
  wire  [31:0] insn_o_2_274_0;
  wire  [31:0] insn_o_2_650_0;
  wire  [31:0] insn_o_2_283_0;
  wire  [31:0] insn_o_2_662_0;
  wire  [31:0] insn_o_2_288_0;
  wire  [31:0] insn_o_2_674_0;
  wire  [31:0] insn_o_2_296_0;
  wire  [31:0] insn_o_2_686_0;
  wire  [31:0] insn_o_2_305_0;
  wire  [31:0] insn_o_2_698_0;
  wire  [31:0] insn_o_2_310_0;
  wire  [31:0] insn_o_2_710_0;
  wire  [31:0] insn_o_2_318_0;
  wire  [31:0] insn_o_2_722_0;
  wire  [31:0] insn_o_2_736_0;
  wire  [31:0] insn_o_2_738_0;
  wire  [31:0] insn_o_2_742_0;
  wire  [31:0] insn_o_2_744_0;
  wire  [31:0] insn_o_2_745_0;
  wire  [31:0] insn_o_2_748_0;
  wire  [31:0] insn_o_2_750_0;
  wire  [31:0] insn_o_2_752_0;
  wire  [16:0] insn_o_2_761_0;
  wire  [14:0] insn_o_2_765_0;
  wire  [31:0] insn_o_2_767_0;
  wire  [31:0] insn_o_2_769_0;
  wire  [18:0] insn_o_2_778_0;
  wire  [12:0] insn_o_2_782_0;
  wire  [31:0] insn_o_2_784_0;
  wire  [31:0] insn_o_2_786_0;
  wire  [31:0] insn_o_2_796_0;
  wire  [31:0] insn_o_2_798_0;
  wire  [31:0] insn_o_2_802_0;
  wire  [31:0] insn_o_2_804_0;
  wire  [31:0] insn_o_2_805_0;
  wire  [31:0] insn_o_2_808_0;
  wire  [31:0] insn_o_2_810_0;
  wire  [31:0] insn_o_2_812_0;
  wire  [6:0] insn_o_2_821_0;
  wire  [24:0] insn_o_2_825_0;
  wire  [31:0] insn_o_2_827_0;
  wire  [31:0] insn_o_2_829_0;
  wire  [17:0] insn_o_2_838_0;
  wire  [13:0] insn_o_2_842_0;
  wire  [31:0] insn_o_2_844_0;
  wire  [31:0] insn_o_2_846_0;
  wire  [31:0] insn_o_2_856_0;
  wire  [31:0] insn_o_2_858_0;
  wire  [31:0] insn_o_2_859_0;
  wire  [31:0] insn_o_2_864_0;
  wire  [31:0] insn_o_2_865_0;
  wire  [31:0] insn_o_2_866_0;
  wire  [31:0] insn_o_2_868_0;
  wire  [31:0] insn_o_2_869_0;
  wire  [31:0] insn_o_2_327_0;
  wire  [31:0] insn_o_2_875_0;
  wire  [31:0] insn_o_2_330_0;
  wire  [31:0] insn_o_2_881_0;
  wire  [31:0] insn_o_2_883_0;
  wire  [31:0] insn_o_2_888_0;
  wire  [31:0] insn_o_2_890_0;
  wire  [31:0] insn_o_2_894_0;
  wire  [31:0] insn_o_2_895_0;
  wire  [31:0] insn_o_2_896_0;
  wire  [31:0] insn_o_2_898_0;
  wire  [31:0] insn_o_2_899_0;
  wire  [31:0] insn_o_2_901_0;
  wire  [31:0] insn_o_2_903_0;
  wire  [31:0] insn_o_2_905_0;
  wire  [31:0] insn_o_2_907_0;
  wire  [31:0] insn_o_2_909_0;
  wire  [31:0] insn_o_2_914_0;
  wire  [31:0] insn_o_2_916_0;
  wire  [31:0] insn_o_2_917_0;
  wire  [31:0] insn_o_2_922_0;
  wire  [31:0] insn_o_2_923_0;
  wire  [31:0] insn_o_2_924_0;
  wire  [31:0] insn_o_2_926_0;
  wire  [31:0] insn_o_2_927_0;
  wire  [31:0] insn_o_2_930_0;
  wire  [31:0] insn_o_2_338_0;
  wire  [31:0] insn_o_2_936_0;
  wire  [31:0] insn_o_2_939_0;
  wire  [31:0] insn_o_2_341_0;
  wire  [31:0] insn_o_2_945_0;
  wire  [31:0] insn_o_2_947_0;
  wire  [31:0] insn_o_2_952_0;
  wire  [31:0] insn_o_2_954_0;
  wire  [31:0] insn_o_2_958_0;
  wire  [31:0] insn_o_2_959_0;
  wire  [31:0] insn_o_2_960_0;
  wire  [31:0] insn_o_2_962_0;
  wire  [31:0] insn_o_2_963_0;
  wire  [31:0] insn_o_2_965_0;
  wire  [31:0] insn_o_2_967_0;
  wire  [31:0] insn_o_2_969_0;
  wire  [31:0] insn_o_2_971_0;
  wire  [31:0] insn_o_2_973_0;
  wire  [31:0] insn_o_2_978_0;
  wire  [31:0] insn_o_2_980_0;
  wire  [31:0] insn_o_2_981_0;
  wire  [31:0] insn_o_2_986_0;
  wire  [31:0] insn_o_2_987_0;
  wire  [31:0] insn_o_2_988_0;
  wire  [31:0] insn_o_2_990_0;
  wire  [31:0] insn_o_2_991_0;
  wire  [31:0] insn_o_2_994_0;
  wire  [31:0] insn_o_2_349_0;
  wire  [31:0] insn_o_2_1000_0;
  wire  [31:0] insn_o_2_1003_0;
  wire  [31:0] insn_o_2_352_0;
  wire  [31:0] insn_o_2_1009_0;
  wire  [31:0] insn_o_2_1011_0;
  wire  [31:0] insn_o_2_1016_0;
  wire  [31:0] insn_o_2_1018_0;
  wire  [31:0] insn_o_2_1022_0;
  wire  [31:0] insn_o_2_1023_0;
  wire  [31:0] insn_o_2_1024_0;
  wire  [31:0] insn_o_2_1026_0;
  wire  [31:0] insn_o_2_1027_0;
  wire  [31:0] insn_o_2_1029_0;
  wire  [31:0] insn_o_2_1031_0;
  wire  [31:0] insn_o_2_1033_0;
  wire  [31:0] insn_o_2_1035_0;
  wire  [31:0] insn_o_2_1037_0;
  wire  [31:0] insn_o_2_1042_0;
  wire  [31:0] insn_o_2_1044_0;
  wire  [31:0] insn_o_2_1045_0;
  wire  [31:0] insn_o_2_1050_0;
  wire  [31:0] insn_o_2_1051_0;
  wire  [31:0] insn_o_2_1052_0;
  wire  [31:0] insn_o_2_1054_0;
  wire  [31:0] insn_o_2_1055_0;
  wire  [31:0] insn_o_2_1058_0;
  wire  [31:0] insn_o_2_360_0;
  wire  [31:0] insn_o_2_1064_0;
  wire  [31:0] insn_o_2_1067_0;
  wire  [31:0] insn_o_2_363_0;
  wire  [31:0] insn_o_2_1073_0;
  wire  [31:0] insn_o_2_1075_0;
  wire  [31:0] insn_o_2_1080_0;
  wire  [31:0] insn_o_2_1082_0;
  wire  [31:0] insn_o_2_1086_0;
  wire  [31:0] insn_o_2_1087_0;
  wire  [31:0] insn_o_2_1088_0;
  wire  [31:0] insn_o_2_1090_0;
  wire  [31:0] insn_o_2_1091_0;
  wire  [31:0] insn_o_2_1093_0;
  wire  [31:0] insn_o_2_1095_0;
  wire  [31:0] insn_o_2_1097_0;
  wire  [31:0] insn_o_2_1099_0;
  wire  [31:0] insn_o_2_1101_0;
  wire  [31:0] insn_o_2_1106_0;
  wire  [31:0] insn_o_2_1108_0;
  wire  [31:0] insn_o_2_1109_0;
  wire  [31:0] insn_o_2_1114_0;
  wire  [31:0] insn_o_2_1115_0;
  wire  [31:0] insn_o_2_1116_0;
  wire  [31:0] insn_o_2_1118_0;
  wire  [31:0] insn_o_2_1119_0;
  wire  [31:0] insn_o_2_1122_0;
  wire  [31:0] insn_o_2_371_0;
  wire  [31:0] insn_o_2_1128_0;
  wire  [31:0] insn_o_2_1131_0;
  wire  [31:0] insn_o_2_374_0;
  wire  [31:0] insn_o_2_1137_0;
  wire  [31:0] insn_o_2_1139_0;
  wire  [31:0] insn_o_2_1144_0;
  wire  [31:0] insn_o_2_1146_0;
  wire  [31:0] insn_o_2_1150_0;
  wire  [31:0] insn_o_2_1151_0;
  wire  [31:0] insn_o_2_1152_0;
  wire  [31:0] insn_o_2_1154_0;
  wire  [31:0] insn_o_2_1155_0;
  wire  [31:0] insn_o_2_1157_0;
  wire  [31:0] insn_o_2_1159_0;
  wire  [31:0] insn_o_2_1161_0;
  wire  [31:0] insn_o_2_1163_0;
  wire  [31:0] insn_o_2_1165_0;
  wire  [31:0] insn_o_2_1170_0;
  wire  [31:0] insn_o_2_1172_0;
  wire  [31:0] insn_o_2_1173_0;
  wire  [31:0] insn_o_2_1178_0;
  wire  [31:0] insn_o_2_1179_0;
  wire  [31:0] insn_o_2_1180_0;
  wire  [31:0] insn_o_2_1182_0;
  wire  [31:0] insn_o_2_1183_0;
  wire  [31:0] insn_o_2_1186_0;
  wire  [31:0] insn_o_2_384_0;
  wire  [31:0] insn_o_2_1192_0;
  wire  [31:0] insn_o_2_1195_0;
  wire  [31:0] insn_o_2_388_0;
  wire  [31:0] insn_o_2_1201_0;
  wire  [31:0] insn_o_2_1203_0;
  wire  [31:0] insn_o_2_1208_0;
  wire  [31:0] insn_o_2_1210_0;
  wire  [31:0] insn_o_2_1214_0;
  wire  [31:0] insn_o_2_1215_0;
  wire  [31:0] insn_o_2_1216_0;
  wire  [31:0] insn_o_2_1218_0;
  wire  [31:0] insn_o_2_1219_0;
  wire  [31:0] insn_o_2_1221_0;
  wire  [31:0] insn_o_2_1223_0;
  wire  [31:0] insn_o_2_1225_0;
  wire  [31:0] insn_o_2_1227_0;
  wire  [31:0] insn_o_2_1229_0;
  wire  [31:0] insn_o_2_1234_0;
  wire  [31:0] insn_o_2_1236_0;
  wire  [31:0] insn_o_2_1237_0;
  wire  [31:0] insn_o_2_1242_0;
  wire  [31:0] insn_o_2_1243_0;
  wire  [31:0] insn_o_2_1244_0;
  wire  [31:0] insn_o_2_1246_0;
  wire  [31:0] insn_o_2_1247_0;
  wire  [31:0] insn_o_2_1250_0;
  wire  [31:0] insn_o_2_391_0;
  wire  [31:0] insn_o_2_1256_0;
  wire  [31:0] insn_o_2_1259_0;
  wire  [31:0] insn_o_2_395_0;
  wire  [31:0] insn_o_2_1265_0;
  wire  [31:0] insn_o_2_1267_0;
  wire  [31:0] insn_o_2_1272_0;
  wire  [31:0] insn_o_2_1274_0;
  wire  [31:0] insn_o_2_1278_0;
  wire  [31:0] insn_o_2_1279_0;
  wire  [31:0] insn_o_2_1280_0;
  wire  [31:0] insn_o_2_1282_0;
  wire  [31:0] insn_o_2_1283_0;
  wire  [31:0] insn_o_2_1285_0;
  wire  [31:0] insn_o_2_1287_0;
  wire  [31:0] insn_o_2_1289_0;
  wire  [31:0] insn_o_2_1291_0;
  wire  [31:0] insn_o_2_1293_0;
  wire  [31:0] insn_o_2_1298_0;
  wire  [31:0] insn_o_2_1300_0;
  wire  [31:0] insn_o_2_1301_0;
  wire  [31:0] insn_o_2_1306_0;
  wire  [31:0] insn_o_2_1307_0;
  wire  [31:0] insn_o_2_1308_0;
  wire  [31:0] insn_o_2_1310_0;
  wire  [31:0] insn_o_2_1311_0;
  wire  [31:0] insn_o_2_1314_0;
  wire  [31:0] insn_o_2_398_0;
  wire  [31:0] insn_o_2_1320_0;
  wire  [31:0] insn_o_2_1323_0;
  wire  [31:0] insn_o_2_402_0;
  wire  [31:0] insn_o_2_1329_0;
  wire  [31:0] insn_o_2_1331_0;
  wire  [31:0] insn_o_2_1336_0;
  wire  [31:0] insn_o_2_1338_0;
  wire  [31:0] insn_o_2_1342_0;
  wire  [31:0] insn_o_2_1343_0;
  wire  [31:0] insn_o_2_1344_0;
  wire  [31:0] insn_o_2_1346_0;
  wire  [31:0] insn_o_2_1347_0;
  wire  [31:0] insn_o_2_1349_0;
  wire  [31:0] insn_o_2_1351_0;
  wire  [31:0] insn_o_2_1353_0;
  wire  [31:0] insn_o_2_1355_0;
  wire  [31:0] insn_o_2_1357_0;
  wire  [31:0] insn_o_2_1359_0;
  wire  [31:0] insn_o_2_1361_0;
  wire  [31:0] insn_o_2_1363_0;
  wire  [31:0] insn_o_2_1365_0;
  wire  [31:0] insn_o_2_1367_0;
  wire  [31:0] insn_o_2_1369_0;
  wire  [31:0] insn_o_2_1371_0;
  wire  [31:0] insn_o_2_1373_0;
  wire  [31:0] insn_o_2_1383_0;
  wire  [31:0] insn_o_2_1385_0;
  wire  [31:0] insn_o_2_1389_0;
  wire  [31:0] insn_o_2_1391_0;
  wire  [31:0] insn_o_2_1392_0;
  wire  [31:0] insn_o_2_1397_0;
  wire  [31:0] insn_o_2_1399_0;
  wire  [31:0] insn_o_2_1400_0;
  wire  [31:0] insn_o_2_1402_0;
  wire  [5:0] insn_o_2_1411_0;
  wire  [25:0] insn_o_2_1415_0;
  wire  [31:0] insn_o_2_1417_0;
  wire  [31:0] insn_o_2_1419_0;
  wire  [10:0] insn_o_2_1428_0;
  wire  [20:0] insn_o_2_1432_0;
  wire  [31:0] insn_o_2_1434_0;
  wire  [31:0] insn_o_2_1436_0;
  wire  [24:0] insn_o_2_1445_0;
  wire  [6:0] insn_o_2_1449_0;
  wire  [31:0] insn_o_2_1451_0;
  wire  [31:0] insn_o_2_1453_0;
  wire  [31:0] insn_o_2_1460_0;
  wire  [31:0] insn_o_2_1462_0;
  wire  [31:0] insn_o_2_1464_0;
  wire  [31:0] insn_o_2_1466_0;
  wire  [31:0] insn_o_2_1476_0;
  wire  [31:0] insn_o_2_1478_0;
  wire  [31:0] insn_o_2_1482_0;
  wire  [31:0] insn_o_2_1484_0;
  wire  [31:0] insn_o_2_1485_0;
  wire  [31:0] insn_o_2_1490_0;
  wire  [31:0] insn_o_2_1492_0;
  wire  [31:0] insn_o_2_1493_0;
  wire  [31:0] insn_o_2_1495_0;
  wire  [1:0] insn_o_2_1504_0;
  wire  [29:0] insn_o_2_1508_0;
  wire  [31:0] insn_o_2_1510_0;
  wire  [31:0] insn_o_2_1512_0;
  wire  [12:0] insn_o_2_1521_0;
  wire  [18:0] insn_o_2_1525_0;
  wire  [31:0] insn_o_2_1527_0;
  wire  [31:0] insn_o_2_1529_0;
  wire  [21:0] insn_o_2_1538_0;
  wire  [9:0] insn_o_2_1542_0;
  wire  [31:0] insn_o_2_1544_0;
  wire  [31:0] insn_o_2_1546_0;
  wire  [31:0] insn_o_2_1553_0;
  wire  [31:0] insn_o_2_1555_0;
  wire  [31:0] insn_o_2_1557_0;
  wire  [31:0] insn_o_2_1559_0;
  wire  [31:0] insn_o_2_1561_0;
  wire  [31:0] insn_o_2_1571_0;
  wire  [31:0] insn_o_2_1573_0;
  wire  [31:0] insn_o_2_1577_0;
  wire  [31:0] insn_o_2_1579_0;
  wire  [31:0] insn_o_2_1580_0;
  wire  [31:0] insn_o_2_1585_0;
  wire  [31:0] insn_o_2_1587_0;
  wire  [31:0] insn_o_2_1588_0;
  wire  [31:0] insn_o_2_1590_0;
  wire  [5:0] insn_o_2_1599_0;
  wire  [25:0] insn_o_2_1603_0;
  wire  [31:0] insn_o_2_1605_0;
  wire  [31:0] insn_o_2_1607_0;
  wire  [10:0] insn_o_2_1616_0;
  wire  [20:0] insn_o_2_1620_0;
  wire  [31:0] insn_o_2_1622_0;
  wire  [31:0] insn_o_2_1624_0;
  wire  [24:0] insn_o_2_1633_0;
  wire  [6:0] insn_o_2_1637_0;
  wire  [31:0] insn_o_2_1639_0;
  wire  [31:0] insn_o_2_1641_0;
  wire  [31:0] insn_o_2_1648_0;
  wire  [31:0] insn_o_2_1650_0;
  wire  [31:0] insn_o_2_1652_0;
  wire  [31:0] insn_o_2_1654_0;
  wire  [31:0] insn_o_2_1664_0;
  wire  [31:0] insn_o_2_1666_0;
  wire  [31:0] insn_o_2_1670_0;
  wire  [31:0] insn_o_2_1672_0;
  wire  [31:0] insn_o_2_1673_0;
  wire  [31:0] insn_o_2_1678_0;
  wire  [31:0] insn_o_2_1680_0;
  wire  [31:0] insn_o_2_1681_0;
  wire  [31:0] insn_o_2_1683_0;
  wire  [1:0] insn_o_2_1692_0;
  wire  [29:0] insn_o_2_1696_0;
  wire  [31:0] insn_o_2_1698_0;
  wire  [31:0] insn_o_2_1700_0;
  wire  [12:0] insn_o_2_1709_0;
  wire  [18:0] insn_o_2_1713_0;
  wire  [31:0] insn_o_2_1715_0;
  wire  [31:0] insn_o_2_1717_0;
  wire  [21:0] insn_o_2_1726_0;
  wire  [9:0] insn_o_2_1730_0;
  wire  [31:0] insn_o_2_1732_0;
  wire  [31:0] insn_o_2_1734_0;
  wire  [31:0] insn_o_2_1741_0;
  wire  [31:0] insn_o_2_1743_0;
  wire  [31:0] insn_o_2_1745_0;
  wire  [31:0] insn_o_2_1747_0;
  wire  [31:0] insn_o_2_1749_0;
  wire  [31:0] insn_o_2_1759_0;
  wire  [31:0] insn_o_2_1761_0;
  wire  [31:0] insn_o_2_1765_0;
  wire  [31:0] insn_o_2_1767_0;
  wire  [31:0] insn_o_2_1768_0;
  wire  [31:0] insn_o_2_1773_0;
  wire  [31:0] insn_o_2_1775_0;
  wire  [31:0] insn_o_2_1776_0;
  wire  [31:0] insn_o_2_1778_0;
  wire  [5:0] insn_o_2_1787_0;
  wire  [25:0] insn_o_2_1791_0;
  wire  [31:0] insn_o_2_1793_0;
  wire  [31:0] insn_o_2_1795_0;
  wire  [10:0] insn_o_2_1804_0;
  wire  [20:0] insn_o_2_1808_0;
  wire  [31:0] insn_o_2_1810_0;
  wire  [31:0] insn_o_2_1812_0;
  wire  [24:0] insn_o_2_1821_0;
  wire  [6:0] insn_o_2_1825_0;
  wire  [31:0] insn_o_2_1827_0;
  wire  [31:0] insn_o_2_1829_0;
  wire  [31:0] insn_o_2_1836_0;
  wire  [31:0] insn_o_2_1838_0;
  wire  [31:0] insn_o_2_1840_0;
  wire  [31:0] insn_o_2_1842_0;
  wire  [31:0] insn_o_2_1852_0;
  wire  [31:0] insn_o_2_1854_0;
  wire  [31:0] insn_o_2_1858_0;
  wire  [31:0] insn_o_2_1860_0;
  wire  [31:0] insn_o_2_1861_0;
  wire  [31:0] insn_o_2_1866_0;
  wire  [31:0] insn_o_2_1868_0;
  wire  [31:0] insn_o_2_1869_0;
  wire  [31:0] insn_o_2_1871_0;
  wire  [1:0] insn_o_2_1880_0;
  wire  [29:0] insn_o_2_1884_0;
  wire  [31:0] insn_o_2_1886_0;
  wire  [31:0] insn_o_2_1888_0;
  wire  [12:0] insn_o_2_1897_0;
  wire  [18:0] insn_o_2_1901_0;
  wire  [31:0] insn_o_2_1903_0;
  wire  [31:0] insn_o_2_1905_0;
  wire  [21:0] insn_o_2_1914_0;
  wire  [9:0] insn_o_2_1918_0;
  wire  [31:0] insn_o_2_1920_0;
  wire  [31:0] insn_o_2_1922_0;
  wire  [31:0] insn_o_2_1929_0;
  wire  [31:0] insn_o_2_1931_0;
  wire  [31:0] insn_o_2_1933_0;
  wire  [31:0] insn_o_2_1935_0;
  wire  [31:0] insn_o_2_1937_0;
  wire  [31:0] insn_o_2_1947_0;
  wire  [31:0] insn_o_2_1949_0;
  wire  [31:0] insn_o_2_1953_0;
  wire  [31:0] insn_o_2_1955_0;
  wire  [31:0] insn_o_2_1956_0;
  wire  [31:0] insn_o_2_1961_0;
  wire  [31:0] insn_o_2_1963_0;
  wire  [31:0] insn_o_2_1964_0;
  wire  [31:0] insn_o_2_1966_0;
  wire  [5:0] insn_o_2_1975_0;
  wire  [25:0] insn_o_2_1979_0;
  wire  [31:0] insn_o_2_1981_0;
  wire  [31:0] insn_o_2_1983_0;
  wire  [10:0] insn_o_2_1992_0;
  wire  [20:0] insn_o_2_1996_0;
  wire  [31:0] insn_o_2_1998_0;
  wire  [31:0] insn_o_2_2000_0;
  wire  [24:0] insn_o_2_2009_0;
  wire  [6:0] insn_o_2_2013_0;
  wire  [31:0] insn_o_2_2015_0;
  wire  [31:0] insn_o_2_2017_0;
  wire  [31:0] insn_o_2_2024_0;
  wire  [31:0] insn_o_2_2026_0;
  wire  [31:0] insn_o_2_2028_0;
  wire  [31:0] insn_o_2_2030_0;
  wire  [31:0] insn_o_2_2040_0;
  wire  [31:0] insn_o_2_2042_0;
  wire  [31:0] insn_o_2_2046_0;
  wire  [31:0] insn_o_2_2048_0;
  wire  [31:0] insn_o_2_2049_0;
  wire  [31:0] insn_o_2_2054_0;
  wire  [31:0] insn_o_2_2056_0;
  wire  [31:0] insn_o_2_2057_0;
  wire  [31:0] insn_o_2_2059_0;
  wire  [1:0] insn_o_2_2068_0;
  wire  [29:0] insn_o_2_2072_0;
  wire  [31:0] insn_o_2_2074_0;
  wire  [31:0] insn_o_2_2076_0;
  wire  [12:0] insn_o_2_2085_0;
  wire  [18:0] insn_o_2_2089_0;
  wire  [31:0] insn_o_2_2091_0;
  wire  [31:0] insn_o_2_2093_0;
  wire  [21:0] insn_o_2_2102_0;
  wire  [9:0] insn_o_2_2106_0;
  wire  [31:0] insn_o_2_2108_0;
  wire  [31:0] insn_o_2_2110_0;
  wire  [31:0] insn_o_2_2117_0;
  wire  [31:0] insn_o_2_2119_0;
  wire  [31:0] insn_o_2_2121_0;
  wire  [31:0] insn_o_2_2123_0;
  wire  [31:0] insn_o_2_2125_0;
  wire  [31:0] insn_o_2_2135_0;
  wire  [31:0] insn_o_2_2137_0;
  wire  [31:0] insn_o_2_2141_0;
  wire  [31:0] insn_o_2_2143_0;
  wire  [31:0] insn_o_2_2144_0;
  wire  [31:0] insn_o_2_2149_0;
  wire  [31:0] insn_o_2_2151_0;
  wire  [31:0] insn_o_2_2152_0;
  wire  [31:0] insn_o_2_2154_0;
  wire  [5:0] insn_o_2_2163_0;
  wire  [25:0] insn_o_2_2167_0;
  wire  [31:0] insn_o_2_2169_0;
  wire  [31:0] insn_o_2_2171_0;
  wire  [10:0] insn_o_2_2180_0;
  wire  [20:0] insn_o_2_2184_0;
  wire  [31:0] insn_o_2_2186_0;
  wire  [31:0] insn_o_2_2188_0;
  wire  [24:0] insn_o_2_2197_0;
  wire  [6:0] insn_o_2_2201_0;
  wire  [31:0] insn_o_2_2203_0;
  wire  [31:0] insn_o_2_2205_0;
  wire  [31:0] insn_o_2_2212_0;
  wire  [31:0] insn_o_2_2214_0;
  wire  [31:0] insn_o_2_2216_0;
  wire  [31:0] insn_o_2_2218_0;
  wire  [31:0] insn_o_2_2228_0;
  wire  [31:0] insn_o_2_2230_0;
  wire  [31:0] insn_o_2_2234_0;
  wire  [31:0] insn_o_2_2236_0;
  wire  [31:0] insn_o_2_2237_0;
  wire  [31:0] insn_o_2_2242_0;
  wire  [31:0] insn_o_2_2244_0;
  wire  [31:0] insn_o_2_2245_0;
  wire  [31:0] insn_o_2_2247_0;
  wire  [1:0] insn_o_2_2256_0;
  wire  [29:0] insn_o_2_2260_0;
  wire  [31:0] insn_o_2_2262_0;
  wire  [31:0] insn_o_2_2264_0;
  wire  [12:0] insn_o_2_2273_0;
  wire  [18:0] insn_o_2_2277_0;
  wire  [31:0] insn_o_2_2279_0;
  wire  [31:0] insn_o_2_2281_0;
  wire  [21:0] insn_o_2_2290_0;
  wire  [9:0] insn_o_2_2294_0;
  wire  [31:0] insn_o_2_2296_0;
  wire  [31:0] insn_o_2_2298_0;
  wire  [31:0] insn_o_2_2305_0;
  wire  [31:0] insn_o_2_2307_0;
  wire  [31:0] insn_o_2_2309_0;
  wire  [31:0] insn_o_2_2311_0;
  wire  [31:0] insn_o_2_2313_0;
  wire  [31:0] insn_o_2_2323_0;
  wire  [31:0] insn_o_2_2325_0;
  wire  [31:0] insn_o_2_2329_0;
  wire  [31:0] insn_o_2_2331_0;
  wire  [31:0] insn_o_2_2332_0;
  wire  [31:0] insn_o_2_2337_0;
  wire  [31:0] insn_o_2_2339_0;
  wire  [31:0] insn_o_2_2340_0;
  wire  [31:0] insn_o_2_2342_0;
  wire  [5:0] insn_o_2_2351_0;
  wire  [25:0] insn_o_2_2355_0;
  wire  [31:0] insn_o_2_2357_0;
  wire  [31:0] insn_o_2_2359_0;
  wire  [10:0] insn_o_2_2368_0;
  wire  [20:0] insn_o_2_2372_0;
  wire  [31:0] insn_o_2_2374_0;
  wire  [31:0] insn_o_2_2376_0;
  wire  [24:0] insn_o_2_2385_0;
  wire  [6:0] insn_o_2_2389_0;
  wire  [31:0] insn_o_2_2391_0;
  wire  [31:0] insn_o_2_2393_0;
  wire  [31:0] insn_o_2_2400_0;
  wire  [31:0] insn_o_2_2402_0;
  wire  [31:0] insn_o_2_2404_0;
  wire  [31:0] insn_o_2_2406_0;
  wire  [31:0] insn_o_2_2416_0;
  wire  [31:0] insn_o_2_2418_0;
  wire  [31:0] insn_o_2_2422_0;
  wire  [31:0] insn_o_2_2424_0;
  wire  [31:0] insn_o_2_2425_0;
  wire  [31:0] insn_o_2_2430_0;
  wire  [31:0] insn_o_2_2432_0;
  wire  [31:0] insn_o_2_2433_0;
  wire  [31:0] insn_o_2_2435_0;
  wire  [1:0] insn_o_2_2444_0;
  wire  [29:0] insn_o_2_2448_0;
  wire  [31:0] insn_o_2_2450_0;
  wire  [31:0] insn_o_2_2452_0;
  wire  [12:0] insn_o_2_2461_0;
  wire  [18:0] insn_o_2_2465_0;
  wire  [31:0] insn_o_2_2467_0;
  wire  [31:0] insn_o_2_2469_0;
  wire  [21:0] insn_o_2_2478_0;
  wire  [9:0] insn_o_2_2482_0;
  wire  [31:0] insn_o_2_2484_0;
  wire  [31:0] insn_o_2_2486_0;
  wire  [31:0] insn_o_2_2493_0;
  wire  [31:0] insn_o_2_2495_0;
  wire  [31:0] insn_o_2_2497_0;
  wire  [31:0] insn_o_2_2499_0;
  wire  [31:0] insn_o_2_2501_0;
  wire  [31:0] insn_o_2_2511_0;
  wire  [31:0] insn_o_2_2513_0;
  wire  [31:0] insn_o_2_2517_0;
  wire  [31:0] insn_o_2_2519_0;
  wire  [31:0] insn_o_2_2520_0;
  wire  [31:0] insn_o_2_2525_0;
  wire  [31:0] insn_o_2_2527_0;
  wire  [31:0] insn_o_2_2528_0;
  wire  [31:0] insn_o_2_2530_0;
  wire  [5:0] insn_o_2_2539_0;
  wire  [25:0] insn_o_2_2543_0;
  wire  [31:0] insn_o_2_2545_0;
  wire  [31:0] insn_o_2_2547_0;
  wire  [10:0] insn_o_2_2556_0;
  wire  [20:0] insn_o_2_2560_0;
  wire  [31:0] insn_o_2_2562_0;
  wire  [31:0] insn_o_2_2564_0;
  wire  [24:0] insn_o_2_2573_0;
  wire  [6:0] insn_o_2_2577_0;
  wire  [31:0] insn_o_2_2579_0;
  wire  [31:0] insn_o_2_2581_0;
  wire  [31:0] insn_o_2_2588_0;
  wire  [31:0] insn_o_2_2590_0;
  wire  [31:0] insn_o_2_2592_0;
  wire  [31:0] insn_o_2_2594_0;
  wire  [31:0] insn_o_2_2604_0;
  wire  [31:0] insn_o_2_2606_0;
  wire  [31:0] insn_o_2_2610_0;
  wire  [31:0] insn_o_2_2612_0;
  wire  [31:0] insn_o_2_2613_0;
  wire  [31:0] insn_o_2_2618_0;
  wire  [31:0] insn_o_2_2620_0;
  wire  [31:0] insn_o_2_2621_0;
  wire  [31:0] insn_o_2_2623_0;
  wire  [1:0] insn_o_2_2632_0;
  wire  [29:0] insn_o_2_2636_0;
  wire  [31:0] insn_o_2_2638_0;
  wire  [31:0] insn_o_2_2640_0;
  wire  [12:0] insn_o_2_2649_0;
  wire  [18:0] insn_o_2_2653_0;
  wire  [31:0] insn_o_2_2655_0;
  wire  [31:0] insn_o_2_2657_0;
  wire  [21:0] insn_o_2_2666_0;
  wire  [9:0] insn_o_2_2670_0;
  wire  [31:0] insn_o_2_2672_0;
  wire  [31:0] insn_o_2_2674_0;
  wire  [31:0] insn_o_2_2681_0;
  wire  [31:0] insn_o_2_2683_0;
  wire  [31:0] insn_o_2_2685_0;
  wire  [31:0] insn_o_2_2687_0;
  wire  [31:0] insn_o_2_2689_0;
  wire  [31:0] insn_o_2_2699_0;
  wire  [31:0] insn_o_2_2701_0;
  wire  [31:0] insn_o_2_2705_0;
  wire  [31:0] insn_o_2_2707_0;
  wire  [31:0] insn_o_2_2708_0;
  wire  [31:0] insn_o_2_2713_0;
  wire  [31:0] insn_o_2_2715_0;
  wire  [31:0] insn_o_2_2716_0;
  wire  [31:0] insn_o_2_2718_0;
  wire  [5:0] insn_o_2_2727_0;
  wire  [25:0] insn_o_2_2731_0;
  wire  [31:0] insn_o_2_2733_0;
  wire  [31:0] insn_o_2_2735_0;
  wire  [10:0] insn_o_2_2744_0;
  wire  [20:0] insn_o_2_2748_0;
  wire  [31:0] insn_o_2_2750_0;
  wire  [31:0] insn_o_2_2752_0;
  wire  [24:0] insn_o_2_2761_0;
  wire  [6:0] insn_o_2_2765_0;
  wire  [31:0] insn_o_2_2767_0;
  wire  [31:0] insn_o_2_2769_0;
  wire  [31:0] insn_o_2_2776_0;
  wire  [31:0] insn_o_2_2778_0;
  wire  [31:0] insn_o_2_2780_0;
  wire  [31:0] insn_o_2_2782_0;
  wire  [31:0] insn_o_2_2792_0;
  wire  [31:0] insn_o_2_2794_0;
  wire  [31:0] insn_o_2_2798_0;
  wire  [31:0] insn_o_2_2800_0;
  wire  [31:0] insn_o_2_2801_0;
  wire  [31:0] insn_o_2_2806_0;
  wire  [31:0] insn_o_2_2808_0;
  wire  [31:0] insn_o_2_2809_0;
  wire  [31:0] insn_o_2_2811_0;
  wire  [1:0] insn_o_2_2820_0;
  wire  [29:0] insn_o_2_2824_0;
  wire  [31:0] insn_o_2_2826_0;
  wire  [31:0] insn_o_2_2828_0;
  wire  [12:0] insn_o_2_2837_0;
  wire  [18:0] insn_o_2_2841_0;
  wire  [31:0] insn_o_2_2843_0;
  wire  [31:0] insn_o_2_2845_0;
  wire  [21:0] insn_o_2_2854_0;
  wire  [9:0] insn_o_2_2858_0;
  wire  [31:0] insn_o_2_2860_0;
  wire  [31:0] insn_o_2_2862_0;
  wire  [31:0] insn_o_2_2869_0;
  wire  [31:0] insn_o_2_2871_0;
  wire  [31:0] insn_o_2_2873_0;
  wire  [31:0] insn_o_2_2875_0;
  wire  [31:0] insn_o_2_2877_0;
  reg [1:0] st_res_2_125;
  reg [1:0] st_res_2_126;
  reg [1:0] st_res_2_193;
  // Insn assigns
  assign insn_o_2_10_0 = gt_124_d0;
  assign insn_o_2_25_0 = add_127_d0;
  assign insn_o_2_29_0 = add_128_d0;
  assign insn_o_2_5_0 = sram_rdata_2;
  assign insn_o_2_39_0 = r50_sha256_237_397[7:0];
  assign insn_o_2_14_0 = sram_rdata_2;
  assign insn_o_2_48_0 = r57_sha256_239_399[15:8];
  assign insn_o_2_50_0 = {r48_sha256_238_398, r55_sha256_240_400};
  assign insn_o_2_19_0 = sram_rdata_2;
  assign insn_o_2_59_0 = r64_sha256_242_402[23:16];
  assign insn_o_2_61_0 = {r47_sha256_241_401, r62_sha256_243_403};
  assign insn_o_2_22_0 = sram_rdata_2;
  assign insn_o_2_70_0 = r71_sha256_245_405[31:24];
  assign insn_o_2_72_0 = {r46_sha256_244_404, r69_sha256_246_406};
  assign insn_o_2_31_0 = sram_rdata_2;
  assign insn_o_2_81_0 = r78_sha256_248_408[7:0];
  assign insn_o_2_83_0 = {r45_sha256_247_407, r76_sha256_249_409};
  assign insn_o_2_35_0 = sram_rdata_2;
  assign insn_o_2_92_0 = r85_sha256_251_411[15:8];
  assign insn_o_2_94_0 = {r44_sha256_250_410, r83_sha256_252_412};
  assign insn_o_2_41_0 = sram_rdata_2;
  assign insn_o_2_103_0 = r92_sha256_254_414[23:16];
  assign insn_o_2_105_0 = {r43_sha256_253_413, r90_sha256_255_415};
  assign insn_o_2_44_0 = sram_rdata_2;
  assign insn_o_2_114_0 = r99_sha256_257_417[31:24];
  assign insn_o_2_116_0 = {r42_sha256_256_416, r97_sha256_258_418};
  assign insn_o_2_52_0 = sram_rdata_2;
  assign insn_o_2_125_0 = r106_sha256_260_420[7:0];
  assign insn_o_2_127_0 = {r41_sha256_259_419, r104_sha256_261_421};
  assign insn_o_2_55_0 = sram_rdata_2;
  assign insn_o_2_136_0 = r113_sha256_263_423[15:8];
  assign insn_o_2_138_0 = {r40_sha256_262_422, r111_sha256_264_424};
  assign insn_o_2_63_0 = sram_rdata_2;
  assign insn_o_2_147_0 = r120_sha256_266_426[23:16];
  assign insn_o_2_149_0 = {r39_sha256_265_425, r118_sha256_267_427};
  assign insn_o_2_66_0 = sram_rdata_2;
  assign insn_o_2_158_0 = r127_sha256_269_429[31:24];
  assign insn_o_2_160_0 = {r38_sha256_268_428, r125_sha256_270_430};
  assign insn_o_2_74_0 = sram_rdata_2;
  assign insn_o_2_169_0 = r134_sha256_272_432[7:0];
  assign insn_o_2_171_0 = {r37_sha256_271_431, r132_sha256_273_433};
  assign insn_o_2_77_0 = sram_rdata_2;
  assign insn_o_2_180_0 = r141_sha256_275_435[15:8];
  assign insn_o_2_182_0 = {r36_sha256_274_434, r139_sha256_276_436};
  assign insn_o_2_85_0 = sram_rdata_2;
  assign insn_o_2_191_0 = r148_sha256_278_438[23:16];
  assign insn_o_2_193_0 = {r35_sha256_277_437, r146_sha256_279_439};
  assign insn_o_2_88_0 = sram_rdata_2;
  assign insn_o_2_202_0 = r155_sha256_281_441[31:24];
  assign insn_o_2_204_0 = {r34_sha256_280_440, r153_sha256_282_442};
  assign insn_o_2_96_0 = sram_rdata_2;
  assign insn_o_2_213_0 = r162_sha256_284_444[7:0];
  assign insn_o_2_215_0 = {r33_sha256_283_443, r160_sha256_285_445};
  assign insn_o_2_99_0 = sram_rdata_2;
  assign insn_o_2_224_0 = r169_sha256_287_447[15:8];
  assign insn_o_2_226_0 = {r32_sha256_286_446, r167_sha256_288_448};
  assign insn_o_2_107_0 = sram_rdata_2;
  assign insn_o_2_235_0 = r176_sha256_290_450[23:16];
  assign insn_o_2_237_0 = {r31_sha256_289_449, r174_sha256_291_451};
  assign insn_o_2_110_0 = sram_rdata_2;
  assign insn_o_2_246_0 = r183_sha256_293_453[31:24];
  assign insn_o_2_248_0 = {r30_sha256_292_452, r181_sha256_294_454};
  assign insn_o_2_118_0 = sram_rdata_2;
  assign insn_o_2_257_0 = r190_sha256_296_456[7:0];
  assign insn_o_2_259_0 = {r29_sha256_295_455, r188_sha256_297_457};
  assign insn_o_2_121_0 = sram_rdata_2;
  assign insn_o_2_268_0 = r197_sha256_299_459[15:8];
  assign insn_o_2_270_0 = {r28_sha256_298_458, r195_sha256_300_460};
  assign insn_o_2_129_0 = sram_rdata_2;
  assign insn_o_2_279_0 = r204_sha256_302_462[23:16];
  assign insn_o_2_281_0 = {r27_sha256_301_461, r202_sha256_303_463};
  assign insn_o_2_132_0 = sram_rdata_2;
  assign insn_o_2_290_0 = r211_sha256_305_465[31:24];
  assign insn_o_2_292_0 = {r26_sha256_304_464, r209_sha256_306_466};
  assign insn_o_2_140_0 = sram_rdata_2;
  assign insn_o_2_301_0 = r218_sha256_308_468[7:0];
  assign insn_o_2_303_0 = {r25_sha256_307_467, r216_sha256_309_469};
  assign insn_o_2_143_0 = sram_rdata_2;
  assign insn_o_2_312_0 = r225_sha256_311_471[15:8];
  assign insn_o_2_314_0 = {r24_sha256_310_470, r223_sha256_312_472};
  assign insn_o_2_151_0 = sram_rdata_2;
  assign insn_o_2_323_0 = r232_sha256_314_474[23:16];
  assign insn_o_2_325_0 = {r23_sha256_313_473, r230_sha256_315_475};
  assign insn_o_2_154_0 = sram_rdata_2;
  assign insn_o_2_334_0 = r239_sha256_317_477[31:24];
  assign insn_o_2_336_0 = {r22_sha256_316_476, r237_sha256_318_478};
  assign insn_o_2_162_0 = sram_rdata_2;
  assign insn_o_2_345_0 = r246_sha256_320_480[7:0];
  assign insn_o_2_347_0 = {r21_sha256_319_479, r244_sha256_321_481};
  assign insn_o_2_165_0 = sram_rdata_2;
  assign insn_o_2_356_0 = r253_sha256_323_483[15:8];
  assign insn_o_2_358_0 = {r20_sha256_322_482, r251_sha256_324_484};
  assign insn_o_2_173_0 = sram_rdata_2;
  assign insn_o_2_367_0 = r260_sha256_326_486[23:16];
  assign insn_o_2_369_0 = {r19_sha256_325_485, r258_sha256_327_487};
  assign insn_o_2_176_0 = sram_rdata_2;
  assign insn_o_2_378_0 = r267_sha256_329_489[31:24];
  assign insn_o_2_380_0 = {r18_sha256_328_488, r265_sha256_330_490};
  assign insn_o_2_445_0 = gt_194_d0;
  assign insn_o_2_450_0 = mem_1_2_125_1_2_125_rbuf;
  assign insn_o_2_456_0 = r1_transform_336_497[7:0];
  assign insn_o_2_460_0 = r1_transform_336_497[15:8];
  assign insn_o_2_462_0 = {r11_transform_337_498, r14_transform_338_499};
  assign insn_o_2_466_0 = r1_transform_336_497[23:16];
  assign insn_o_2_468_0 = {r10_transform_339_500, r17_transform_340_501};
  assign insn_o_2_472_0 = r1_transform_336_497[31:24];
  assign insn_o_2_474_0 = {r9_transform_341_502, r20_transform_342_503};
  assign insn_o_2_480_0 = add_202_d0;
  assign insn_o_2_487_0 = gt_203_d0;
  assign insn_o_2_492_0 = sub_204_d0;
  assign insn_o_2_198_0 = sram_rdata_223;
  assign insn_o_2_504_0 = sub_205_d0;
  assign insn_o_2_206_0 = sram_rdata_223;
  assign insn_o_2_510_0 = add_206_d0;
  assign insn_o_2_514_0 = sub_207_d0;
  assign insn_o_2_209_0 = sram_rdata_223;
  assign insn_o_2_525_0 = add_208_d0;
  assign insn_o_2_528_0 = sub_209_d0;
  assign insn_o_2_217_0 = sram_rdata_223;
  assign insn_o_2_534_0 = add_210_d0;
  assign insn_o_2_540_0 = add_211_d0;
  assign insn_o_2_222_0 = sram_rdata_2;
  assign insn_o_2_229_0 = sram_rdata_2;
  assign insn_o_2_233_0 = sram_rdata_2;
  assign insn_o_2_240_0 = sram_rdata_2;
  assign insn_o_2_244_0 = sram_rdata_2;
  assign insn_o_2_251_0 = sram_rdata_2;
  assign insn_o_2_255_0 = sram_rdata_2;
  assign insn_o_2_262_0 = sram_rdata_2;
  assign insn_o_2_603_0 = gt_212_d0;
  assign insn_o_2_628_0 = add_213_d0;
  assign insn_o_2_266_0 = sram_rdata_2;
  assign insn_o_2_638_0 = add_214_d0;
  assign insn_o_2_274_0 = sram_rdata_2;
  assign insn_o_2_650_0 = add_215_d0;
  assign insn_o_2_283_0 = sram_rdata_2;
  assign insn_o_2_662_0 = add_216_d0;
  assign insn_o_2_288_0 = sram_rdata_2;
  assign insn_o_2_674_0 = add_217_d0;
  assign insn_o_2_296_0 = sram_rdata_2;
  assign insn_o_2_686_0 = add_218_d0;
  assign insn_o_2_305_0 = sram_rdata_2;
  assign insn_o_2_698_0 = add_219_d0;
  assign insn_o_2_310_0 = sram_rdata_2;
  assign insn_o_2_710_0 = add_220_d0;
  assign insn_o_2_318_0 = sram_rdata_2;
  assign insn_o_2_722_0 = add_221_d0;
  assign insn_o_2_745_0 = r4_s1_226_555 ^ r6_s1_227_556;
  assign insn_o_2_748_0 = x_224_554 >> 10;
  assign insn_o_2_750_0 = r3_s1_228_557 ^ r8_s1_229_558;
  assign insn_o_2_761_0 = arg_177_561[16:0];
  assign insn_o_2_765_0 = arg_177_561[31:17];
  assign insn_o_2_767_0 = {r3_ror32_17_179_562, r6_ror32_17_180_563};
  assign insn_o_2_778_0 = arg_187_566[18:0];
  assign insn_o_2_782_0 = arg_187_566[31:19];
  assign insn_o_2_784_0 = {r3_ror32_19_189_567, r6_ror32_19_190_568};
  assign insn_o_2_805_0 = r4_s0_219_572 ^ r6_s0_220_573;
  assign insn_o_2_808_0 = x_217_571 >> 3;
  assign insn_o_2_810_0 = r3_s0_221_574 ^ r8_s0_222_575;
  assign insn_o_2_821_0 = arg_212_578[6:0];
  assign insn_o_2_825_0 = arg_212_578[31:7];
  assign insn_o_2_827_0 = {r3_ror32_7_214_579, r6_ror32_7_215_580};
  assign insn_o_2_838_0 = arg_182_583[17:0];
  assign insn_o_2_842_0 = arg_182_583[31:18];
  assign insn_o_2_844_0 = {r3_ror32_18_184_584, r6_ror32_18_185_585};
  assign insn_o_2_859_0 = add_16_d0;
  assign insn_o_2_869_0 = add_17_d0;
  assign insn_o_2_327_0 = sram_rdata_222;
  assign insn_o_2_875_0 = add_19_d0;
  assign insn_o_2_330_0 = sram_rdata_223;
  assign insn_o_2_881_0 = add_21_d0;
  assign insn_o_2_899_0 = add_22_d0;
  assign insn_o_2_903_0 = add_23_d0;
  assign insn_o_2_907_0 = add_24_d0;
  assign insn_o_2_917_0 = add_25_d0;
  assign insn_o_2_927_0 = add_26_d0;
  assign insn_o_2_930_0 = add_27_d0;
  assign insn_o_2_338_0 = sram_rdata_222;
  assign insn_o_2_936_0 = add_28_d0;
  assign insn_o_2_939_0 = add_29_d0;
  assign insn_o_2_341_0 = sram_rdata_223;
  assign insn_o_2_945_0 = add_30_d0;
  assign insn_o_2_963_0 = add_31_d0;
  assign insn_o_2_967_0 = add_32_d0;
  assign insn_o_2_971_0 = add_33_d0;
  assign insn_o_2_981_0 = add_34_d0;
  assign insn_o_2_991_0 = add_35_d0;
  assign insn_o_2_994_0 = add_36_d0;
  assign insn_o_2_349_0 = sram_rdata_222;
  assign insn_o_2_1000_0 = add_37_d0;
  assign insn_o_2_1003_0 = add_38_d0;
  assign insn_o_2_352_0 = sram_rdata_223;
  assign insn_o_2_1009_0 = add_39_d0;
  assign insn_o_2_1027_0 = add_40_d0;
  assign insn_o_2_1031_0 = add_41_d0;
  assign insn_o_2_1035_0 = add_42_d0;
  assign insn_o_2_1045_0 = add_43_d0;
  assign insn_o_2_1055_0 = add_44_d0;
  assign insn_o_2_1058_0 = add_45_d0;
  assign insn_o_2_360_0 = sram_rdata_222;
  assign insn_o_2_1064_0 = add_46_d0;
  assign insn_o_2_1067_0 = add_47_d0;
  assign insn_o_2_363_0 = sram_rdata_223;
  assign insn_o_2_1073_0 = add_48_d0;
  assign insn_o_2_1091_0 = add_49_d0;
  assign insn_o_2_1095_0 = add_50_d0;
  assign insn_o_2_1099_0 = add_51_d0;
  assign insn_o_2_1109_0 = add_52_d0;
  assign insn_o_2_1119_0 = add_53_d0;
  assign insn_o_2_1122_0 = add_54_d0;
  assign insn_o_2_371_0 = sram_rdata_222;
  assign insn_o_2_1128_0 = add_55_d0;
  assign insn_o_2_1131_0 = add_56_d0;
  assign insn_o_2_374_0 = sram_rdata_223;
  assign insn_o_2_1137_0 = add_57_d0;
  assign insn_o_2_1155_0 = add_58_d0;
  assign insn_o_2_1159_0 = add_59_d0;
  assign insn_o_2_1163_0 = add_60_d0;
  assign insn_o_2_1173_0 = add_61_d0;
  assign insn_o_2_1183_0 = add_62_d0;
  assign insn_o_2_1186_0 = add_63_d0;
  assign insn_o_2_384_0 = sram_rdata_222;
  assign insn_o_2_1192_0 = add_64_d0;
  assign insn_o_2_1195_0 = add_65_d0;
  assign insn_o_2_388_0 = sram_rdata_223;
  assign insn_o_2_1201_0 = add_66_d0;
  assign insn_o_2_1219_0 = add_67_d0;
  assign insn_o_2_1223_0 = add_68_d0;
  assign insn_o_2_1227_0 = add_69_d0;
  assign insn_o_2_1237_0 = add_70_d0;
  assign insn_o_2_1247_0 = add_71_d0;
  assign insn_o_2_1250_0 = add_72_d0;
  assign insn_o_2_391_0 = sram_rdata_222;
  assign insn_o_2_1256_0 = add_73_d0;
  assign insn_o_2_1259_0 = add_74_d0;
  assign insn_o_2_395_0 = sram_rdata_223;
  assign insn_o_2_1265_0 = add_75_d0;
  assign insn_o_2_1283_0 = add_76_d0;
  assign insn_o_2_1287_0 = add_77_d0;
  assign insn_o_2_1291_0 = add_78_d0;
  assign insn_o_2_1301_0 = add_79_d0;
  assign insn_o_2_1311_0 = add_80_d0;
  assign insn_o_2_1314_0 = add_81_d0;
  assign insn_o_2_398_0 = sram_rdata_222;
  assign insn_o_2_1320_0 = add_82_d0;
  assign insn_o_2_1323_0 = add_83_d0;
  assign insn_o_2_402_0 = sram_rdata_223;
  assign insn_o_2_1329_0 = add_84_d0;
  assign insn_o_2_1347_0 = add_85_d0;
  assign insn_o_2_1351_0 = add_86_d0;
  assign insn_o_2_1355_0 = add_87_d0;
  assign insn_o_2_1392_0 = r4_e1_24_726 ^ r6_e1_25_727;
  assign insn_o_2_1400_0 = r3_e1_26_728 ^ r8_e1_27_729;
  assign insn_o_2_1411_0 = arg_207_732[5:0];
  assign insn_o_2_1415_0 = arg_207_732[31:6];
  assign insn_o_2_1417_0 = {r3_ror32_6_209_733, r6_ror32_6_210_734};
  assign insn_o_2_1428_0 = arg_167_737[10:0];
  assign insn_o_2_1432_0 = arg_167_737[31:11];
  assign insn_o_2_1434_0 = {r3_ror32_11_169_738, r6_ror32_11_170_739};
  assign insn_o_2_1445_0 = arg_202_742[24:0];
  assign insn_o_2_1449_0 = arg_202_742[31:25];
  assign insn_o_2_1451_0 = {r3_ror32_25_204_743, r6_ror32_25_205_744};
  assign insn_o_2_1460_0 = y_1_747 ^ z_2_748;
  assign insn_o_2_1462_0 = x_0_750 & r6_Ch_4_749;
  assign insn_o_2_1464_0 = z_2_748 ^ r5_Ch_5_751;
  assign insn_o_2_1485_0 = r4_e0_17_755 ^ r6_e0_18_756;
  assign insn_o_2_1493_0 = r3_e0_19_757 ^ r8_e0_20_758;
  assign insn_o_2_1504_0 = arg_192_761[1:0];
  assign insn_o_2_1508_0 = arg_192_761[31:2];
  assign insn_o_2_1510_0 = {r3_ror32_2_194_762, r6_ror32_2_195_763};
  assign insn_o_2_1521_0 = arg_172_766[12:0];
  assign insn_o_2_1525_0 = arg_172_766[31:13];
  assign insn_o_2_1527_0 = {r3_ror32_13_174_767, r6_ror32_13_175_768};
  assign insn_o_2_1538_0 = arg_197_771[21:0];
  assign insn_o_2_1542_0 = arg_197_771[31:22];
  assign insn_o_2_1544_0 = {r3_ror32_22_199_772, r6_ror32_22_200_773};
  assign insn_o_2_1553_0 = x_7_776 & y_8_777;
  assign insn_o_2_1555_0 = x_7_776 | y_8_777;
  assign insn_o_2_1557_0 = z_9_780 & r7_Maj_12_779;
  assign insn_o_2_1559_0 = r5_Maj_11_778 | r6_Maj_13_781;
  assign insn_o_2_1580_0 = r4_e1_24_785 ^ r6_e1_25_786;
  assign insn_o_2_1588_0 = r3_e1_26_787 ^ r8_e1_27_788;
  assign insn_o_2_1599_0 = arg_207_791[5:0];
  assign insn_o_2_1603_0 = arg_207_791[31:6];
  assign insn_o_2_1605_0 = {r3_ror32_6_209_792, r6_ror32_6_210_793};
  assign insn_o_2_1616_0 = arg_167_796[10:0];
  assign insn_o_2_1620_0 = arg_167_796[31:11];
  assign insn_o_2_1622_0 = {r3_ror32_11_169_797, r6_ror32_11_170_798};
  assign insn_o_2_1633_0 = arg_202_801[24:0];
  assign insn_o_2_1637_0 = arg_202_801[31:25];
  assign insn_o_2_1639_0 = {r3_ror32_25_204_802, r6_ror32_25_205_803};
  assign insn_o_2_1648_0 = y_1_806 ^ z_2_807;
  assign insn_o_2_1650_0 = x_0_809 & r6_Ch_4_808;
  assign insn_o_2_1652_0 = z_2_807 ^ r5_Ch_5_810;
  assign insn_o_2_1673_0 = r4_e0_17_814 ^ r6_e0_18_815;
  assign insn_o_2_1681_0 = r3_e0_19_816 ^ r8_e0_20_817;
  assign insn_o_2_1692_0 = arg_192_820[1:0];
  assign insn_o_2_1696_0 = arg_192_820[31:2];
  assign insn_o_2_1698_0 = {r3_ror32_2_194_821, r6_ror32_2_195_822};
  assign insn_o_2_1709_0 = arg_172_825[12:0];
  assign insn_o_2_1713_0 = arg_172_825[31:13];
  assign insn_o_2_1715_0 = {r3_ror32_13_174_826, r6_ror32_13_175_827};
  assign insn_o_2_1726_0 = arg_197_830[21:0];
  assign insn_o_2_1730_0 = arg_197_830[31:22];
  assign insn_o_2_1732_0 = {r3_ror32_22_199_831, r6_ror32_22_200_832};
  assign insn_o_2_1741_0 = x_7_835 & y_8_836;
  assign insn_o_2_1743_0 = x_7_835 | y_8_836;
  assign insn_o_2_1745_0 = z_9_839 & r7_Maj_12_838;
  assign insn_o_2_1747_0 = r5_Maj_11_837 | r6_Maj_13_840;
  assign insn_o_2_1768_0 = r4_e1_24_844 ^ r6_e1_25_845;
  assign insn_o_2_1776_0 = r3_e1_26_846 ^ r8_e1_27_847;
  assign insn_o_2_1787_0 = arg_207_850[5:0];
  assign insn_o_2_1791_0 = arg_207_850[31:6];
  assign insn_o_2_1793_0 = {r3_ror32_6_209_851, r6_ror32_6_210_852};
  assign insn_o_2_1804_0 = arg_167_855[10:0];
  assign insn_o_2_1808_0 = arg_167_855[31:11];
  assign insn_o_2_1810_0 = {r3_ror32_11_169_856, r6_ror32_11_170_857};
  assign insn_o_2_1821_0 = arg_202_860[24:0];
  assign insn_o_2_1825_0 = arg_202_860[31:25];
  assign insn_o_2_1827_0 = {r3_ror32_25_204_861, r6_ror32_25_205_862};
  assign insn_o_2_1836_0 = y_1_865 ^ z_2_866;
  assign insn_o_2_1838_0 = x_0_868 & r6_Ch_4_867;
  assign insn_o_2_1840_0 = z_2_866 ^ r5_Ch_5_869;
  assign insn_o_2_1861_0 = r4_e0_17_873 ^ r6_e0_18_874;
  assign insn_o_2_1869_0 = r3_e0_19_875 ^ r8_e0_20_876;
  assign insn_o_2_1880_0 = arg_192_879[1:0];
  assign insn_o_2_1884_0 = arg_192_879[31:2];
  assign insn_o_2_1886_0 = {r3_ror32_2_194_880, r6_ror32_2_195_881};
  assign insn_o_2_1897_0 = arg_172_884[12:0];
  assign insn_o_2_1901_0 = arg_172_884[31:13];
  assign insn_o_2_1903_0 = {r3_ror32_13_174_885, r6_ror32_13_175_886};
  assign insn_o_2_1914_0 = arg_197_889[21:0];
  assign insn_o_2_1918_0 = arg_197_889[31:22];
  assign insn_o_2_1920_0 = {r3_ror32_22_199_890, r6_ror32_22_200_891};
  assign insn_o_2_1929_0 = x_7_894 & y_8_895;
  assign insn_o_2_1931_0 = x_7_894 | y_8_895;
  assign insn_o_2_1933_0 = z_9_898 & r7_Maj_12_897;
  assign insn_o_2_1935_0 = r5_Maj_11_896 | r6_Maj_13_899;
  assign insn_o_2_1956_0 = r4_e1_24_903 ^ r6_e1_25_904;
  assign insn_o_2_1964_0 = r3_e1_26_905 ^ r8_e1_27_906;
  assign insn_o_2_1975_0 = arg_207_909[5:0];
  assign insn_o_2_1979_0 = arg_207_909[31:6];
  assign insn_o_2_1981_0 = {r3_ror32_6_209_910, r6_ror32_6_210_911};
  assign insn_o_2_1992_0 = arg_167_914[10:0];
  assign insn_o_2_1996_0 = arg_167_914[31:11];
  assign insn_o_2_1998_0 = {r3_ror32_11_169_915, r6_ror32_11_170_916};
  assign insn_o_2_2009_0 = arg_202_919[24:0];
  assign insn_o_2_2013_0 = arg_202_919[31:25];
  assign insn_o_2_2015_0 = {r3_ror32_25_204_920, r6_ror32_25_205_921};
  assign insn_o_2_2024_0 = y_1_924 ^ z_2_925;
  assign insn_o_2_2026_0 = x_0_927 & r6_Ch_4_926;
  assign insn_o_2_2028_0 = z_2_925 ^ r5_Ch_5_928;
  assign insn_o_2_2049_0 = r4_e0_17_932 ^ r6_e0_18_933;
  assign insn_o_2_2057_0 = r3_e0_19_934 ^ r8_e0_20_935;
  assign insn_o_2_2068_0 = arg_192_938[1:0];
  assign insn_o_2_2072_0 = arg_192_938[31:2];
  assign insn_o_2_2074_0 = {r3_ror32_2_194_939, r6_ror32_2_195_940};
  assign insn_o_2_2085_0 = arg_172_943[12:0];
  assign insn_o_2_2089_0 = arg_172_943[31:13];
  assign insn_o_2_2091_0 = {r3_ror32_13_174_944, r6_ror32_13_175_945};
  assign insn_o_2_2102_0 = arg_197_948[21:0];
  assign insn_o_2_2106_0 = arg_197_948[31:22];
  assign insn_o_2_2108_0 = {r3_ror32_22_199_949, r6_ror32_22_200_950};
  assign insn_o_2_2117_0 = x_7_953 & y_8_954;
  assign insn_o_2_2119_0 = x_7_953 | y_8_954;
  assign insn_o_2_2121_0 = z_9_957 & r7_Maj_12_956;
  assign insn_o_2_2123_0 = r5_Maj_11_955 | r6_Maj_13_958;
  assign insn_o_2_2144_0 = r4_e1_24_962 ^ r6_e1_25_963;
  assign insn_o_2_2152_0 = r3_e1_26_964 ^ r8_e1_27_965;
  assign insn_o_2_2163_0 = arg_207_968[5:0];
  assign insn_o_2_2167_0 = arg_207_968[31:6];
  assign insn_o_2_2169_0 = {r3_ror32_6_209_969, r6_ror32_6_210_970};
  assign insn_o_2_2180_0 = arg_167_973[10:0];
  assign insn_o_2_2184_0 = arg_167_973[31:11];
  assign insn_o_2_2186_0 = {r3_ror32_11_169_974, r6_ror32_11_170_975};
  assign insn_o_2_2197_0 = arg_202_978[24:0];
  assign insn_o_2_2201_0 = arg_202_978[31:25];
  assign insn_o_2_2203_0 = {r3_ror32_25_204_979, r6_ror32_25_205_980};
  assign insn_o_2_2212_0 = y_1_983 ^ z_2_984;
  assign insn_o_2_2214_0 = x_0_986 & r6_Ch_4_985;
  assign insn_o_2_2216_0 = z_2_984 ^ r5_Ch_5_987;
  assign insn_o_2_2237_0 = r4_e0_17_991 ^ r6_e0_18_992;
  assign insn_o_2_2245_0 = r3_e0_19_993 ^ r8_e0_20_994;
  assign insn_o_2_2256_0 = arg_192_997[1:0];
  assign insn_o_2_2260_0 = arg_192_997[31:2];
  assign insn_o_2_2262_0 = {r3_ror32_2_194_998, r6_ror32_2_195_999};
  assign insn_o_2_2273_0 = arg_172_1002[12:0];
  assign insn_o_2_2277_0 = arg_172_1002[31:13];
  assign insn_o_2_2279_0 = {r3_ror32_13_174_1003, r6_ror32_13_175_1004};
  assign insn_o_2_2290_0 = arg_197_1007[21:0];
  assign insn_o_2_2294_0 = arg_197_1007[31:22];
  assign insn_o_2_2296_0 = {r3_ror32_22_199_1008, r6_ror32_22_200_1009};
  assign insn_o_2_2305_0 = x_7_1012 & y_8_1013;
  assign insn_o_2_2307_0 = x_7_1012 | y_8_1013;
  assign insn_o_2_2309_0 = z_9_1016 & r7_Maj_12_1015;
  assign insn_o_2_2311_0 = r5_Maj_11_1014 | r6_Maj_13_1017;
  assign insn_o_2_2332_0 = r4_e1_24_1021 ^ r6_e1_25_1022;
  assign insn_o_2_2340_0 = r3_e1_26_1023 ^ r8_e1_27_1024;
  assign insn_o_2_2351_0 = arg_207_1027[5:0];
  assign insn_o_2_2355_0 = arg_207_1027[31:6];
  assign insn_o_2_2357_0 = {r3_ror32_6_209_1028, r6_ror32_6_210_1029};
  assign insn_o_2_2368_0 = arg_167_1032[10:0];
  assign insn_o_2_2372_0 = arg_167_1032[31:11];
  assign insn_o_2_2374_0 = {r3_ror32_11_169_1033, r6_ror32_11_170_1034};
  assign insn_o_2_2385_0 = arg_202_1037[24:0];
  assign insn_o_2_2389_0 = arg_202_1037[31:25];
  assign insn_o_2_2391_0 = {r3_ror32_25_204_1038, r6_ror32_25_205_1039};
  assign insn_o_2_2400_0 = y_1_1042 ^ z_2_1043;
  assign insn_o_2_2402_0 = x_0_1045 & r6_Ch_4_1044;
  assign insn_o_2_2404_0 = z_2_1043 ^ r5_Ch_5_1046;
  assign insn_o_2_2425_0 = r4_e0_17_1050 ^ r6_e0_18_1051;
  assign insn_o_2_2433_0 = r3_e0_19_1052 ^ r8_e0_20_1053;
  assign insn_o_2_2444_0 = arg_192_1056[1:0];
  assign insn_o_2_2448_0 = arg_192_1056[31:2];
  assign insn_o_2_2450_0 = {r3_ror32_2_194_1057, r6_ror32_2_195_1058};
  assign insn_o_2_2461_0 = arg_172_1061[12:0];
  assign insn_o_2_2465_0 = arg_172_1061[31:13];
  assign insn_o_2_2467_0 = {r3_ror32_13_174_1062, r6_ror32_13_175_1063};
  assign insn_o_2_2478_0 = arg_197_1066[21:0];
  assign insn_o_2_2482_0 = arg_197_1066[31:22];
  assign insn_o_2_2484_0 = {r3_ror32_22_199_1067, r6_ror32_22_200_1068};
  assign insn_o_2_2493_0 = x_7_1071 & y_8_1072;
  assign insn_o_2_2495_0 = x_7_1071 | y_8_1072;
  assign insn_o_2_2497_0 = z_9_1075 & r7_Maj_12_1074;
  assign insn_o_2_2499_0 = r5_Maj_11_1073 | r6_Maj_13_1076;
  assign insn_o_2_2520_0 = r4_e1_24_1080 ^ r6_e1_25_1081;
  assign insn_o_2_2528_0 = r3_e1_26_1082 ^ r8_e1_27_1083;
  assign insn_o_2_2539_0 = arg_207_1086[5:0];
  assign insn_o_2_2543_0 = arg_207_1086[31:6];
  assign insn_o_2_2545_0 = {r3_ror32_6_209_1087, r6_ror32_6_210_1088};
  assign insn_o_2_2556_0 = arg_167_1091[10:0];
  assign insn_o_2_2560_0 = arg_167_1091[31:11];
  assign insn_o_2_2562_0 = {r3_ror32_11_169_1092, r6_ror32_11_170_1093};
  assign insn_o_2_2573_0 = arg_202_1096[24:0];
  assign insn_o_2_2577_0 = arg_202_1096[31:25];
  assign insn_o_2_2579_0 = {r3_ror32_25_204_1097, r6_ror32_25_205_1098};
  assign insn_o_2_2588_0 = y_1_1101 ^ z_2_1102;
  assign insn_o_2_2590_0 = x_0_1104 & r6_Ch_4_1103;
  assign insn_o_2_2592_0 = z_2_1102 ^ r5_Ch_5_1105;
  assign insn_o_2_2613_0 = r4_e0_17_1109 ^ r6_e0_18_1110;
  assign insn_o_2_2621_0 = r3_e0_19_1111 ^ r8_e0_20_1112;
  assign insn_o_2_2632_0 = arg_192_1115[1:0];
  assign insn_o_2_2636_0 = arg_192_1115[31:2];
  assign insn_o_2_2638_0 = {r3_ror32_2_194_1116, r6_ror32_2_195_1117};
  assign insn_o_2_2649_0 = arg_172_1120[12:0];
  assign insn_o_2_2653_0 = arg_172_1120[31:13];
  assign insn_o_2_2655_0 = {r3_ror32_13_174_1121, r6_ror32_13_175_1122};
  assign insn_o_2_2666_0 = arg_197_1125[21:0];
  assign insn_o_2_2670_0 = arg_197_1125[31:22];
  assign insn_o_2_2672_0 = {r3_ror32_22_199_1126, r6_ror32_22_200_1127};
  assign insn_o_2_2681_0 = x_7_1130 & y_8_1131;
  assign insn_o_2_2683_0 = x_7_1130 | y_8_1131;
  assign insn_o_2_2685_0 = z_9_1134 & r7_Maj_12_1133;
  assign insn_o_2_2687_0 = r5_Maj_11_1132 | r6_Maj_13_1135;
  assign insn_o_2_2708_0 = r4_e1_24_1139 ^ r6_e1_25_1140;
  assign insn_o_2_2716_0 = r3_e1_26_1141 ^ r8_e1_27_1142;
  assign insn_o_2_2727_0 = arg_207_1145[5:0];
  assign insn_o_2_2731_0 = arg_207_1145[31:6];
  assign insn_o_2_2733_0 = {r3_ror32_6_209_1146, r6_ror32_6_210_1147};
  assign insn_o_2_2744_0 = arg_167_1150[10:0];
  assign insn_o_2_2748_0 = arg_167_1150[31:11];
  assign insn_o_2_2750_0 = {r3_ror32_11_169_1151, r6_ror32_11_170_1152};
  assign insn_o_2_2761_0 = arg_202_1155[24:0];
  assign insn_o_2_2765_0 = arg_202_1155[31:25];
  assign insn_o_2_2767_0 = {r3_ror32_25_204_1156, r6_ror32_25_205_1157};
  assign insn_o_2_2776_0 = y_1_1160 ^ z_2_1161;
  assign insn_o_2_2778_0 = x_0_1163 & r6_Ch_4_1162;
  assign insn_o_2_2780_0 = z_2_1161 ^ r5_Ch_5_1164;
  assign insn_o_2_2801_0 = r4_e0_17_1168 ^ r6_e0_18_1169;
  assign insn_o_2_2809_0 = r3_e0_19_1170 ^ r8_e0_20_1171;
  assign insn_o_2_2820_0 = arg_192_1174[1:0];
  assign insn_o_2_2824_0 = arg_192_1174[31:2];
  assign insn_o_2_2826_0 = {r3_ror32_2_194_1175, r6_ror32_2_195_1176};
  assign insn_o_2_2837_0 = arg_172_1179[12:0];
  assign insn_o_2_2841_0 = arg_172_1179[31:13];
  assign insn_o_2_2843_0 = {r3_ror32_13_174_1180, r6_ror32_13_175_1181};
  assign insn_o_2_2854_0 = arg_197_1184[21:0];
  assign insn_o_2_2858_0 = arg_197_1184[31:22];
  assign insn_o_2_2860_0 = {r3_ror32_22_199_1185, r6_ror32_22_200_1186};
  assign insn_o_2_2869_0 = x_7_1189 & y_8_1190;
  assign insn_o_2_2871_0 = x_7_1189 | y_8_1190;
  assign insn_o_2_2873_0 = z_9_1193 & r7_Maj_12_1192;
  assign insn_o_2_2875_0 = r5_Maj_11_1191 | r6_Maj_13_1194;
  assign insn_o_2_2_0 = ext_task_arg_2_0;
  assign insn_o_2_2_1 = ext_task_arg_2_1;

  // Table 1
  always @(posedge clk) begin
    if (rst) begin
      st_1 <= `S_1_1;
    end else begin
      case (st_1)
        `S_1_1: begin
          st_1 <= `S_1_2;
        end
        `S_1_2: begin
        end
      endcase
    end
  end
  // Table 2
  always @(posedge clk) begin
    if (rst) begin
      st_2 <= `S_2_task_idle;
      mem_1_2_125_1_2_125_ack <= 0;
      mem_1_2_125_1_2_125_req <= 0;
      mem_1_2_125_1_2_125_p0_wen <= 0;
      axi_addr2_126 <= 0;
      axi_wen2_126 <= 0;
      axi_req2_126 <= 0;
      sha256_req_ready <= 0;
      sha256_res_valid <= 0;
      sha256_req_busy <= 0;
      st_res_2_125 <= 0;
      st_res_2_126 <= 0;
      st_res_2_193 <= 0;
    end else begin
      mem_1_2_125_1_2_125_ack <= !(0) && mem_1_2_125_1_2_125_req;
      mem_1_2_125_1_2_125_req <= ((st_2 == `S_2_335 && st_res_2_125 == 0)) && !mem_1_2_125_1_2_125_ack;
      mem_1_2_125_1_2_125_p0_wen <= 0 && !mem_1_2_125_1_2_125_ack;
      axi_req2_126 <= ((st_2 == `S_2_13 && st_res_2_126 == 0)) && !axi_ack2_126;
      axi_wen2_126 <= 0;
      sha256_req_ready <= sha256_req_valid & (st_2 == `S_2_task_idle);
      sha256_req_busy <= !(st_2 == `S_2_task_idle);
      sram_wdata_en_2 <= (st_2 == 519) | (st_2 == 288) | (st_2 == 293) | (st_2 == 298) | (st_2 == 303) | (st_2 == 308) | (st_2 == 313) | (st_2 == 318) | (st_2 == 323) | (st_2 == 456) | (st_2 == 465) | (st_2 == 474) | (st_2 == 483) | (st_2 == 492) | (st_2 == 501) | (st_2 == 510);
      sram_wdata_en_222 <= 0;
      sram_wdata_en_223 <= (st_2 == 354) | (st_2 == 393);
      case (st_2)
        `S_2_task_idle: begin
          if (sha256_req_valid) begin
            st_2 <= `S_2_1;
            ext_task_arg_2_0 <= sha256_req_0;
            ext_task_arg_2_1 <= sha256_req_1;
          end
        end
        `S_2_1: begin
          addr_231_392 <= insn_o_2_2_0;
          blocks_232_393 <= insn_o_2_2_1;
          st_2 <= `S_2_288;
        end
        `S_2_6: begin
          r5_sha256_234_394 <= 32'd0;
          st_2 <= `S_2_7;
        end
        `S_2_7: begin
          r7_sha256_235_395 <= insn_o_2_10_0;
          st_2 <= `S_2_8;
        end
        `S_2_8: begin
          if (r7_sha256_235_395) begin
            st_2 <= `S_2_9;
          end else begin
            st_2 <= `S_2_23;
          end
        end
        `S_2_9: begin
          st_2 <= `S_2_13;
        end
        `S_2_13: begin
          // AXI access request
          if (st_res_2_126 == 0) begin
            axi_addr2_126 <= addr_231_392;
            axi_len2_126 <= 32'd15;
            axi_start2_126 <= 32'd0;
            if (axi_ack2_126) begin
              st_res_2_126 <= 3;
            end
          end
          if ((st_res_2_126 == 3)) begin
            // 1 cycle insns
          end
          if ((st_res_2_126 == 3)) begin
            // clears sub states
            st_res_2_126 <= 0;
          end
          if ((st_res_2_126 == 3)) begin
          st_2 <= `S_2_329;
          end
        end
        `S_2_19: begin
          r16_sha256_236_396 <= insn_o_2_25_0;
          st_2 <= `S_2_20;
        end
        `S_2_20: begin
          addr_231_392 <= r16_sha256_236_396;
          st_2 <= `S_2_21;
        end
        `S_2_21: begin
          r5_sha256_234_394 <= insn_o_2_29_0;
          st_2 <= `S_2_7;
        end
        `S_2_23: begin
          st_2 <= `S_2_26;
        end
        `S_2_26: begin
          sram_addr_2 <= 32'd7;
          st_2 <= `S_2_2;
        end
        `S_2_2: begin
          r50_sha256_237_397 <= insn_o_2_5_0;
          st_2 <= `S_2_29;
        end
        `S_2_29: begin
          r48_sha256_238_398 <= insn_o_2_39_0;
          st_2 <= `S_2_33;
        end
        `S_2_33: begin
          sram_addr_2 <= 32'd7;
          st_2 <= `S_2_3;
        end
        `S_2_3: begin
          r57_sha256_239_399 <= insn_o_2_14_0;
          st_2 <= `S_2_36;
        end
        `S_2_36: begin
          r55_sha256_240_400 <= insn_o_2_48_0;
          st_2 <= `S_2_37;
        end
        `S_2_37: begin
          r47_sha256_241_401 <= insn_o_2_50_0;
          st_2 <= `S_2_41;
        end
        `S_2_41: begin
          sram_addr_2 <= 32'd7;
          st_2 <= `S_2_4;
        end
        `S_2_4: begin
          r64_sha256_242_402 <= insn_o_2_19_0;
          st_2 <= `S_2_44;
        end
        `S_2_44: begin
          r62_sha256_243_403 <= insn_o_2_59_0;
          st_2 <= `S_2_45;
        end
        `S_2_45: begin
          r46_sha256_244_404 <= insn_o_2_61_0;
          st_2 <= `S_2_49;
        end
        `S_2_49: begin
          sram_addr_2 <= 32'd7;
          st_2 <= `S_2_5;
        end
        `S_2_5: begin
          r71_sha256_245_405 <= insn_o_2_22_0;
          st_2 <= `S_2_52;
        end
        `S_2_52: begin
          r69_sha256_246_406 <= insn_o_2_70_0;
          st_2 <= `S_2_53;
        end
        `S_2_53: begin
          r45_sha256_247_407 <= insn_o_2_72_0;
          st_2 <= `S_2_57;
        end
        `S_2_57: begin
          sram_addr_2 <= 32'd6;
          st_2 <= `S_2_10;
        end
        `S_2_10: begin
          r78_sha256_248_408 <= insn_o_2_31_0;
          st_2 <= `S_2_60;
        end
        `S_2_60: begin
          r76_sha256_249_409 <= insn_o_2_81_0;
          st_2 <= `S_2_61;
        end
        `S_2_61: begin
          r44_sha256_250_410 <= insn_o_2_83_0;
          st_2 <= `S_2_65;
        end
        `S_2_65: begin
          sram_addr_2 <= 32'd6;
          st_2 <= `S_2_11;
        end
        `S_2_11: begin
          r85_sha256_251_411 <= insn_o_2_35_0;
          st_2 <= `S_2_68;
        end
        `S_2_68: begin
          r83_sha256_252_412 <= insn_o_2_92_0;
          st_2 <= `S_2_69;
        end
        `S_2_69: begin
          r43_sha256_253_413 <= insn_o_2_94_0;
          st_2 <= `S_2_73;
        end
        `S_2_73: begin
          sram_addr_2 <= 32'd6;
          st_2 <= `S_2_12;
        end
        `S_2_12: begin
          r92_sha256_254_414 <= insn_o_2_41_0;
          st_2 <= `S_2_76;
        end
        `S_2_76: begin
          r90_sha256_255_415 <= insn_o_2_103_0;
          st_2 <= `S_2_77;
        end
        `S_2_77: begin
          r42_sha256_256_416 <= insn_o_2_105_0;
          st_2 <= `S_2_81;
        end
        `S_2_81: begin
          sram_addr_2 <= 32'd6;
          st_2 <= `S_2_14;
        end
        `S_2_14: begin
          r99_sha256_257_417 <= insn_o_2_44_0;
          st_2 <= `S_2_84;
        end
        `S_2_84: begin
          r97_sha256_258_418 <= insn_o_2_114_0;
          st_2 <= `S_2_85;
        end
        `S_2_85: begin
          r41_sha256_259_419 <= insn_o_2_116_0;
          st_2 <= `S_2_89;
        end
        `S_2_89: begin
          sram_addr_2 <= 32'd5;
          st_2 <= `S_2_15;
        end
        `S_2_15: begin
          r106_sha256_260_420 <= insn_o_2_52_0;
          st_2 <= `S_2_92;
        end
        `S_2_92: begin
          r104_sha256_261_421 <= insn_o_2_125_0;
          st_2 <= `S_2_93;
        end
        `S_2_93: begin
          r40_sha256_262_422 <= insn_o_2_127_0;
          st_2 <= `S_2_97;
        end
        `S_2_97: begin
          sram_addr_2 <= 32'd5;
          st_2 <= `S_2_16;
        end
        `S_2_16: begin
          r113_sha256_263_423 <= insn_o_2_55_0;
          st_2 <= `S_2_100;
        end
        `S_2_100: begin
          r111_sha256_264_424 <= insn_o_2_136_0;
          st_2 <= `S_2_101;
        end
        `S_2_101: begin
          r39_sha256_265_425 <= insn_o_2_138_0;
          st_2 <= `S_2_105;
        end
        `S_2_105: begin
          sram_addr_2 <= 32'd5;
          st_2 <= `S_2_17;
        end
        `S_2_17: begin
          r120_sha256_266_426 <= insn_o_2_63_0;
          st_2 <= `S_2_108;
        end
        `S_2_108: begin
          r118_sha256_267_427 <= insn_o_2_147_0;
          st_2 <= `S_2_109;
        end
        `S_2_109: begin
          r38_sha256_268_428 <= insn_o_2_149_0;
          st_2 <= `S_2_113;
        end
        `S_2_113: begin
          sram_addr_2 <= 32'd5;
          st_2 <= `S_2_18;
        end
        `S_2_18: begin
          r127_sha256_269_429 <= insn_o_2_66_0;
          st_2 <= `S_2_116;
        end
        `S_2_116: begin
          r125_sha256_270_430 <= insn_o_2_158_0;
          st_2 <= `S_2_117;
        end
        `S_2_117: begin
          r37_sha256_271_431 <= insn_o_2_160_0;
          st_2 <= `S_2_121;
        end
        `S_2_121: begin
          sram_addr_2 <= 32'd4;
          st_2 <= `S_2_22;
        end
        `S_2_22: begin
          r134_sha256_272_432 <= insn_o_2_74_0;
          st_2 <= `S_2_124;
        end
        `S_2_124: begin
          r132_sha256_273_433 <= insn_o_2_169_0;
          st_2 <= `S_2_125;
        end
        `S_2_125: begin
          r36_sha256_274_434 <= insn_o_2_171_0;
          st_2 <= `S_2_129;
        end
        `S_2_129: begin
          sram_addr_2 <= 32'd4;
          st_2 <= `S_2_24;
        end
        `S_2_24: begin
          r141_sha256_275_435 <= insn_o_2_77_0;
          st_2 <= `S_2_132;
        end
        `S_2_132: begin
          r139_sha256_276_436 <= insn_o_2_180_0;
          st_2 <= `S_2_133;
        end
        `S_2_133: begin
          r35_sha256_277_437 <= insn_o_2_182_0;
          st_2 <= `S_2_137;
        end
        `S_2_137: begin
          sram_addr_2 <= 32'd4;
          st_2 <= `S_2_25;
        end
        `S_2_25: begin
          r148_sha256_278_438 <= insn_o_2_85_0;
          st_2 <= `S_2_140;
        end
        `S_2_140: begin
          r146_sha256_279_439 <= insn_o_2_191_0;
          st_2 <= `S_2_141;
        end
        `S_2_141: begin
          r34_sha256_280_440 <= insn_o_2_193_0;
          st_2 <= `S_2_145;
        end
        `S_2_145: begin
          sram_addr_2 <= 32'd4;
          st_2 <= `S_2_27;
        end
        `S_2_27: begin
          r155_sha256_281_441 <= insn_o_2_88_0;
          st_2 <= `S_2_148;
        end
        `S_2_148: begin
          r153_sha256_282_442 <= insn_o_2_202_0;
          st_2 <= `S_2_149;
        end
        `S_2_149: begin
          r33_sha256_283_443 <= insn_o_2_204_0;
          st_2 <= `S_2_153;
        end
        `S_2_153: begin
          sram_addr_2 <= 32'd3;
          st_2 <= `S_2_28;
        end
        `S_2_28: begin
          r162_sha256_284_444 <= insn_o_2_96_0;
          st_2 <= `S_2_156;
        end
        `S_2_156: begin
          r160_sha256_285_445 <= insn_o_2_213_0;
          st_2 <= `S_2_157;
        end
        `S_2_157: begin
          r32_sha256_286_446 <= insn_o_2_215_0;
          st_2 <= `S_2_161;
        end
        `S_2_161: begin
          sram_addr_2 <= 32'd3;
          st_2 <= `S_2_30;
        end
        `S_2_30: begin
          r169_sha256_287_447 <= insn_o_2_99_0;
          st_2 <= `S_2_164;
        end
        `S_2_164: begin
          r167_sha256_288_448 <= insn_o_2_224_0;
          st_2 <= `S_2_165;
        end
        `S_2_165: begin
          r31_sha256_289_449 <= insn_o_2_226_0;
          st_2 <= `S_2_169;
        end
        `S_2_169: begin
          sram_addr_2 <= 32'd3;
          st_2 <= `S_2_31;
        end
        `S_2_31: begin
          r176_sha256_290_450 <= insn_o_2_107_0;
          st_2 <= `S_2_172;
        end
        `S_2_172: begin
          r174_sha256_291_451 <= insn_o_2_235_0;
          st_2 <= `S_2_173;
        end
        `S_2_173: begin
          r30_sha256_292_452 <= insn_o_2_237_0;
          st_2 <= `S_2_177;
        end
        `S_2_177: begin
          sram_addr_2 <= 32'd3;
          st_2 <= `S_2_32;
        end
        `S_2_32: begin
          r183_sha256_293_453 <= insn_o_2_110_0;
          st_2 <= `S_2_180;
        end
        `S_2_180: begin
          r181_sha256_294_454 <= insn_o_2_246_0;
          st_2 <= `S_2_181;
        end
        `S_2_181: begin
          r29_sha256_295_455 <= insn_o_2_248_0;
          st_2 <= `S_2_185;
        end
        `S_2_185: begin
          sram_addr_2 <= 32'd2;
          st_2 <= `S_2_34;
        end
        `S_2_34: begin
          r190_sha256_296_456 <= insn_o_2_118_0;
          st_2 <= `S_2_188;
        end
        `S_2_188: begin
          r188_sha256_297_457 <= insn_o_2_257_0;
          st_2 <= `S_2_189;
        end
        `S_2_189: begin
          r28_sha256_298_458 <= insn_o_2_259_0;
          st_2 <= `S_2_193;
        end
        `S_2_193: begin
          sram_addr_2 <= 32'd2;
          st_2 <= `S_2_35;
        end
        `S_2_35: begin
          r197_sha256_299_459 <= insn_o_2_121_0;
          st_2 <= `S_2_196;
        end
        `S_2_196: begin
          r195_sha256_300_460 <= insn_o_2_268_0;
          st_2 <= `S_2_197;
        end
        `S_2_197: begin
          r27_sha256_301_461 <= insn_o_2_270_0;
          st_2 <= `S_2_201;
        end
        `S_2_201: begin
          sram_addr_2 <= 32'd2;
          st_2 <= `S_2_38;
        end
        `S_2_38: begin
          r204_sha256_302_462 <= insn_o_2_129_0;
          st_2 <= `S_2_204;
        end
        `S_2_204: begin
          r202_sha256_303_463 <= insn_o_2_279_0;
          st_2 <= `S_2_205;
        end
        `S_2_205: begin
          r26_sha256_304_464 <= insn_o_2_281_0;
          st_2 <= `S_2_209;
        end
        `S_2_209: begin
          sram_addr_2 <= 32'd2;
          st_2 <= `S_2_39;
        end
        `S_2_39: begin
          r211_sha256_305_465 <= insn_o_2_132_0;
          st_2 <= `S_2_212;
        end
        `S_2_212: begin
          r209_sha256_306_466 <= insn_o_2_290_0;
          st_2 <= `S_2_213;
        end
        `S_2_213: begin
          r25_sha256_307_467 <= insn_o_2_292_0;
          st_2 <= `S_2_217;
        end
        `S_2_217: begin
          sram_addr_2 <= 32'd1;
          st_2 <= `S_2_40;
        end
        `S_2_40: begin
          r218_sha256_308_468 <= insn_o_2_140_0;
          st_2 <= `S_2_220;
        end
        `S_2_220: begin
          r216_sha256_309_469 <= insn_o_2_301_0;
          st_2 <= `S_2_221;
        end
        `S_2_221: begin
          r24_sha256_310_470 <= insn_o_2_303_0;
          st_2 <= `S_2_225;
        end
        `S_2_225: begin
          sram_addr_2 <= 32'd1;
          st_2 <= `S_2_42;
        end
        `S_2_42: begin
          r225_sha256_311_471 <= insn_o_2_143_0;
          st_2 <= `S_2_228;
        end
        `S_2_228: begin
          r223_sha256_312_472 <= insn_o_2_312_0;
          st_2 <= `S_2_229;
        end
        `S_2_229: begin
          r23_sha256_313_473 <= insn_o_2_314_0;
          st_2 <= `S_2_233;
        end
        `S_2_233: begin
          sram_addr_2 <= 32'd1;
          st_2 <= `S_2_43;
        end
        `S_2_43: begin
          r232_sha256_314_474 <= insn_o_2_151_0;
          st_2 <= `S_2_236;
        end
        `S_2_236: begin
          r230_sha256_315_475 <= insn_o_2_323_0;
          st_2 <= `S_2_237;
        end
        `S_2_237: begin
          r22_sha256_316_476 <= insn_o_2_325_0;
          st_2 <= `S_2_241;
        end
        `S_2_241: begin
          sram_addr_2 <= 32'd1;
          st_2 <= `S_2_46;
        end
        `S_2_46: begin
          r239_sha256_317_477 <= insn_o_2_154_0;
          st_2 <= `S_2_244;
        end
        `S_2_244: begin
          r237_sha256_318_478 <= insn_o_2_334_0;
          st_2 <= `S_2_245;
        end
        `S_2_245: begin
          r21_sha256_319_479 <= insn_o_2_336_0;
          st_2 <= `S_2_249;
        end
        `S_2_249: begin
          sram_addr_2 <= 32'd0;
          st_2 <= `S_2_47;
        end
        `S_2_47: begin
          r246_sha256_320_480 <= insn_o_2_162_0;
          st_2 <= `S_2_252;
        end
        `S_2_252: begin
          r244_sha256_321_481 <= insn_o_2_345_0;
          st_2 <= `S_2_253;
        end
        `S_2_253: begin
          r20_sha256_322_482 <= insn_o_2_347_0;
          st_2 <= `S_2_257;
        end
        `S_2_257: begin
          sram_addr_2 <= 32'd0;
          st_2 <= `S_2_48;
        end
        `S_2_48: begin
          r253_sha256_323_483 <= insn_o_2_165_0;
          st_2 <= `S_2_260;
        end
        `S_2_260: begin
          r251_sha256_324_484 <= insn_o_2_356_0;
          st_2 <= `S_2_261;
        end
        `S_2_261: begin
          r19_sha256_325_485 <= insn_o_2_358_0;
          st_2 <= `S_2_265;
        end
        `S_2_265: begin
          sram_addr_2 <= 32'd0;
          st_2 <= `S_2_50;
        end
        `S_2_50: begin
          r260_sha256_326_486 <= insn_o_2_173_0;
          st_2 <= `S_2_268;
        end
        `S_2_268: begin
          r258_sha256_327_487 <= insn_o_2_367_0;
          st_2 <= `S_2_269;
        end
        `S_2_269: begin
          r18_sha256_328_488 <= insn_o_2_369_0;
          st_2 <= `S_2_273;
        end
        `S_2_273: begin
          sram_addr_2 <= 32'd0;
          st_2 <= `S_2_51;
        end
        `S_2_51: begin
          r267_sha256_329_489 <= insn_o_2_176_0;
          st_2 <= `S_2_276;
        end
        `S_2_276: begin
          r265_sha256_330_490 <= insn_o_2_378_0;
          st_2 <= `S_2_277;
        end
        `S_2_277: begin
          r17_sha256_331_491 <= insn_o_2_380_0;
          st_2 <= `S_2_278;
        end
        `S_2_278: begin
          r2_sha256_233_492 <= r17_sha256_331_491;
          st_2 <= `S_2_282;
        end
        `S_2_282: begin
          if (st_res_2_193 == 0) begin
            sha256_res_valid <= 1;
            st_res_2_193 <= 1;
            sha256_res_0 <= r2_sha256_233_492;
          end
          if (st_res_2_193 == 1) begin
            if (sha256_res_ready) begin
              sha256_res_valid <= 0;
              st_res_2_193 <= 3;
            end
          end
          if ((st_res_2_193 == 3)) begin
            // 1 cycle insns
          end
          if ((st_res_2_193 == 3)) begin
            // clears sub states
            st_res_2_193 <= 0;
          end
          if ((st_res_2_193 == 3)) begin
          st_2 <= `S_2_task_idle;
          end
        end
        `S_2_288: begin
          sram_addr_2 <= 32'd0;
          sram_wdata_2 <= 32'd1779033703;
          st_2 <= `S_2_293;
        end
        `S_2_293: begin
          sram_addr_2 <= 32'd1;
          sram_wdata_2 <= 32'd2147483647;
          st_2 <= `S_2_298;
        end
        `S_2_298: begin
          sram_addr_2 <= 32'd2;
          sram_wdata_2 <= 32'd1013904242;
          st_2 <= `S_2_303;
        end
        `S_2_303: begin
          sram_addr_2 <= 32'd3;
          sram_wdata_2 <= 32'd2147483647;
          st_2 <= `S_2_308;
        end
        `S_2_308: begin
          sram_addr_2 <= 32'd4;
          sram_wdata_2 <= 32'd1359893119;
          st_2 <= `S_2_313;
        end
        `S_2_313: begin
          sram_addr_2 <= 32'd5;
          sram_wdata_2 <= 32'd2147483647;
          st_2 <= `S_2_318;
        end
        `S_2_318: begin
          sram_addr_2 <= 32'd6;
          sram_wdata_2 <= 32'd528734635;
          st_2 <= `S_2_323;
        end
        `S_2_323: begin
          sram_addr_2 <= 32'd7;
          sram_wdata_2 <= 32'd1541459225;
          st_2 <= `S_2_6;
        end
        `S_2_329: begin
          r0_transform_333_494 <= 32'd0;
          st_2 <= `S_2_330;
        end
        `S_2_330: begin
          st_2 <= `S_2_331;
        end
        `S_2_331: begin
          r3_transform_334_495 <= insn_o_2_445_0;
          st_2 <= `S_2_332;
        end
        `S_2_332: begin
          if (r3_transform_334_495) begin
            st_2 <= `S_2_333;
          end else begin
            st_2 <= `S_2_357;
          end
        end
        `S_2_333: begin
          st_2 <= `S_2_335;
        end
        `S_2_335: begin
          if (st_res_2_125 == 0) begin
            mem_1_2_125_1_2_125_p0_addr <= r0_transform_333_494;
            if (mem_1_2_125_1_2_125_ack) begin
              st_res_2_125 <= 3;
              mem_1_2_125_1_2_125_rbuf <= mem_1_2_125_p0_rdata;
            end
          end
          if ((st_res_2_125 == 3)) begin
            // 1 cycle insns
          r5_transform_335_496 <= insn_o_2_450_0;
          end
          if ((st_res_2_125 == 3)) begin
            // clears sub states
            st_res_2_125 <= 0;
          end
          if ((st_res_2_125 == 3)) begin
          st_2 <= `S_2_336;
          end
        end
        `S_2_336: begin
          r1_transform_336_497 <= r5_transform_335_496;
          st_2 <= `S_2_339;
        end
        `S_2_339: begin
          r11_transform_337_498 <= insn_o_2_456_0;
          st_2 <= `S_2_342;
        end
        `S_2_342: begin
          r14_transform_338_499 <= insn_o_2_460_0;
          st_2 <= `S_2_343;
        end
        `S_2_343: begin
          r10_transform_339_500 <= insn_o_2_462_0;
          st_2 <= `S_2_346;
        end
        `S_2_346: begin
          r17_transform_340_501 <= insn_o_2_466_0;
          st_2 <= `S_2_347;
        end
        `S_2_347: begin
          r9_transform_341_502 <= insn_o_2_468_0;
          st_2 <= `S_2_350;
        end
        `S_2_350: begin
          r20_transform_342_503 <= insn_o_2_472_0;
          st_2 <= `S_2_351;
        end
        `S_2_351: begin
          r8_transform_343_504 <= insn_o_2_474_0;
          st_2 <= `S_2_354;
        end
        `S_2_354: begin
          sram_addr_223 <= r0_transform_333_494;
          sram_wdata_223 <= r8_transform_343_504;
          st_2 <= `S_2_355;
        end
        `S_2_355: begin
          r0_transform_333_494 <= insn_o_2_480_0;
          st_2 <= `S_2_330;
        end
        `S_2_357: begin
          st_2 <= `S_2_358;
        end
        `S_2_358: begin
          r0_transform_333_494 <= 32'd16;
          st_2 <= `S_2_359;
        end
        `S_2_359: begin
          st_2 <= `S_2_360;
        end
        `S_2_360: begin
          r26_transform_344_505 <= insn_o_2_487_0;
          st_2 <= `S_2_361;
        end
        `S_2_361: begin
          if (r26_transform_344_505) begin
            st_2 <= `S_2_362;
          end else begin
            st_2 <= `S_2_396;
          end
        end
        `S_2_362: begin
          st_2 <= `S_2_364;
        end
        `S_2_364: begin
          r33_transform_345_506 <= insn_o_2_492_0;
          st_2 <= `S_2_367;
        end
        `S_2_367: begin
          sram_addr_223 <= r33_transform_345_506;
          st_2 <= `S_2_54;
        end
        `S_2_54: begin
          r35_transform_346_507 <= insn_o_2_198_0;
          st_2 <= `S_2_368;
        end
        `S_2_368: begin
          x_224_554 <= r35_transform_346_507;
          st_2 <= `S_2_525;
        end
        `S_2_369: begin
          r31_transform_347_508 <= r1_s1_225_560;
          st_2 <= `S_2_371;
        end
        `S_2_371: begin
          r38_transform_348_509 <= insn_o_2_504_0;
          st_2 <= `S_2_374;
        end
        `S_2_374: begin
          sram_addr_223 <= r38_transform_348_509;
          st_2 <= `S_2_55;
        end
        `S_2_55: begin
          r40_transform_349_510 <= insn_o_2_206_0;
          st_2 <= `S_2_375;
        end
        `S_2_375: begin
          r30_transform_350_511 <= insn_o_2_510_0;
          st_2 <= `S_2_378;
        end
        `S_2_378: begin
          r45_transform_351_512 <= insn_o_2_514_0;
          st_2 <= `S_2_381;
        end
        `S_2_381: begin
          sram_addr_223 <= r45_transform_351_512;
          st_2 <= `S_2_56;
        end
        `S_2_56: begin
          r47_transform_352_513 <= insn_o_2_209_0;
          st_2 <= `S_2_382;
        end
        `S_2_382: begin
          x_217_571 <= r47_transform_352_513;
          st_2 <= `S_2_567;
        end
        `S_2_383: begin
          r43_transform_353_514 <= r1_s0_218_577;
          st_2 <= `S_2_384;
        end
        `S_2_384: begin
          r29_transform_354_515 <= insn_o_2_525_0;
          st_2 <= `S_2_386;
        end
        `S_2_386: begin
          r50_transform_355_516 <= insn_o_2_528_0;
          st_2 <= `S_2_389;
        end
        `S_2_389: begin
          sram_addr_223 <= r50_transform_355_516;
          st_2 <= `S_2_58;
        end
        `S_2_58: begin
          r52_transform_356_517 <= insn_o_2_217_0;
          st_2 <= `S_2_390;
        end
        `S_2_390: begin
          r28_transform_357_518 <= insn_o_2_534_0;
          st_2 <= `S_2_393;
        end
        `S_2_393: begin
          sram_addr_223 <= r0_transform_333_494;
          sram_wdata_223 <= r28_transform_357_518;
          st_2 <= `S_2_394;
        end
        `S_2_394: begin
          r0_transform_333_494 <= insn_o_2_540_0;
          st_2 <= `S_2_359;
        end
        `S_2_396: begin
          st_2 <= `S_2_399;
        end
        `S_2_399: begin
          sram_addr_2 <= 32'd0;
          st_2 <= `S_2_59;
        end
        `S_2_59: begin
          r66_transform_358_519 <= insn_o_2_222_0;
          st_2 <= `S_2_400;
        end
        `S_2_400: begin
          r57_transform_359_520 <= r66_transform_358_519;
          st_2 <= `S_2_404;
        end
        `S_2_404: begin
          sram_addr_2 <= 32'd1;
          st_2 <= `S_2_62;
        end
        `S_2_62: begin
          r70_transform_360_521 <= insn_o_2_229_0;
          st_2 <= `S_2_405;
        end
        `S_2_405: begin
          r58_transform_361_522 <= r70_transform_360_521;
          st_2 <= `S_2_409;
        end
        `S_2_409: begin
          sram_addr_2 <= 32'd2;
          st_2 <= `S_2_63;
        end
        `S_2_63: begin
          r74_transform_362_523 <= insn_o_2_233_0;
          st_2 <= `S_2_410;
        end
        `S_2_410: begin
          r59_transform_363_524 <= r74_transform_362_523;
          st_2 <= `S_2_414;
        end
        `S_2_414: begin
          sram_addr_2 <= 32'd3;
          st_2 <= `S_2_64;
        end
        `S_2_64: begin
          r78_transform_364_525 <= insn_o_2_240_0;
          st_2 <= `S_2_415;
        end
        `S_2_415: begin
          r60_transform_365_526 <= r78_transform_364_525;
          st_2 <= `S_2_419;
        end
        `S_2_419: begin
          sram_addr_2 <= 32'd4;
          st_2 <= `S_2_66;
        end
        `S_2_66: begin
          r82_transform_366_527 <= insn_o_2_244_0;
          st_2 <= `S_2_420;
        end
        `S_2_420: begin
          r61_transform_367_528 <= r82_transform_366_527;
          st_2 <= `S_2_424;
        end
        `S_2_424: begin
          sram_addr_2 <= 32'd5;
          st_2 <= `S_2_67;
        end
        `S_2_67: begin
          r86_transform_368_529 <= insn_o_2_251_0;
          st_2 <= `S_2_425;
        end
        `S_2_425: begin
          r62_transform_369_530 <= r86_transform_368_529;
          st_2 <= `S_2_429;
        end
        `S_2_429: begin
          sram_addr_2 <= 32'd6;
          st_2 <= `S_2_70;
        end
        `S_2_70: begin
          r90_transform_370_531 <= insn_o_2_255_0;
          st_2 <= `S_2_430;
        end
        `S_2_430: begin
          r63_transform_371_532 <= r90_transform_370_531;
          st_2 <= `S_2_434;
        end
        `S_2_434: begin
          sram_addr_2 <= 32'd7;
          st_2 <= `S_2_71;
        end
        `S_2_71: begin
          r94_transform_372_533 <= insn_o_2_262_0;
          st_2 <= `S_2_435;
        end
        `S_2_435: begin
          r64_transform_373_534 <= r94_transform_372_533;
          st_2 <= `S_2_437;
        end
        `S_2_437: begin
          r0_transform_333_494 <= 32'd0;
          st_2 <= `S_2_438;
        end
        `S_2_438: begin
          st_2 <= `S_2_439;
        end
        `S_2_439: begin
          r98_transform_374_535 <= insn_o_2_603_0;
          st_2 <= `S_2_440;
        end
        `S_2_440: begin
          if (r98_transform_374_535) begin
            st_2 <= `S_2_441;
          end else begin
            st_2 <= `S_2_448;
          end
        end
        `S_2_441: begin
          st_2 <= `S_2_442;
        end
        `S_2_442: begin
          a_30_602 <= r57_transform_359_520;
          b_31_604 <= r58_transform_361_522;
          c_32_605 <= r59_transform_363_524;
          d_33_609 <= r60_transform_365_526;
          e_34_588 <= r61_transform_367_528;
          f_35_592 <= r62_transform_369_530;
          g_36_593 <= r63_transform_371_532;
          h_37_590 <= r64_transform_373_534;
          idx_38_596 <= r0_transform_333_494;
          st_2 <= `S_2_609;
        end
        `S_2_443: begin
          r57_transform_359_520 <= r9_iterate_39_717;
          r58_transform_361_522 <= r10_iterate_40_718;
          r59_transform_363_524 <= r11_iterate_41_719;
          r60_transform_365_526 <= r12_iterate_42_720;
          r61_transform_367_528 <= r13_iterate_43_721;
          r62_transform_369_530 <= r14_iterate_44_722;
          r63_transform_371_532 <= r15_iterate_45_723;
          r64_transform_373_534 <= r16_iterate_46_724;
          st_2 <= `S_2_445;
        end
        `S_2_445: begin
          r102_transform_375_536 <= insn_o_2_628_0;
          st_2 <= `S_2_446;
        end
        `S_2_446: begin
          r0_transform_333_494 <= r102_transform_375_536;
          st_2 <= `S_2_438;
        end
        `S_2_448: begin
          st_2 <= `S_2_451;
        end
        `S_2_451: begin
          sram_addr_2 <= 32'd0;
          st_2 <= `S_2_72;
        end
        `S_2_72: begin
          r104_transform_376_537 <= insn_o_2_266_0;
          st_2 <= `S_2_452;
        end
        `S_2_452: begin
          r107_transform_377_538 <= insn_o_2_638_0;
          st_2 <= `S_2_456;
        end
        `S_2_456: begin
          sram_addr_2 <= 32'd0;
          sram_wdata_2 <= r107_transform_377_538;
          st_2 <= `S_2_460;
        end
        `S_2_460: begin
          sram_addr_2 <= 32'd1;
          st_2 <= `S_2_74;
        end
        `S_2_74: begin
          r112_transform_378_539 <= insn_o_2_274_0;
          st_2 <= `S_2_461;
        end
        `S_2_461: begin
          r115_transform_379_540 <= insn_o_2_650_0;
          st_2 <= `S_2_465;
        end
        `S_2_465: begin
          sram_addr_2 <= 32'd1;
          sram_wdata_2 <= r115_transform_379_540;
          st_2 <= `S_2_469;
        end
        `S_2_469: begin
          sram_addr_2 <= 32'd2;
          st_2 <= `S_2_75;
        end
        `S_2_75: begin
          r120_transform_380_541 <= insn_o_2_283_0;
          st_2 <= `S_2_470;
        end
        `S_2_470: begin
          r123_transform_381_542 <= insn_o_2_662_0;
          st_2 <= `S_2_474;
        end
        `S_2_474: begin
          sram_addr_2 <= 32'd2;
          sram_wdata_2 <= r123_transform_381_542;
          st_2 <= `S_2_478;
        end
        `S_2_478: begin
          sram_addr_2 <= 32'd3;
          st_2 <= `S_2_78;
        end
        `S_2_78: begin
          r128_transform_382_543 <= insn_o_2_288_0;
          st_2 <= `S_2_479;
        end
        `S_2_479: begin
          r131_transform_383_544 <= insn_o_2_674_0;
          st_2 <= `S_2_483;
        end
        `S_2_483: begin
          sram_addr_2 <= 32'd3;
          sram_wdata_2 <= r131_transform_383_544;
          st_2 <= `S_2_487;
        end
        `S_2_487: begin
          sram_addr_2 <= 32'd4;
          st_2 <= `S_2_79;
        end
        `S_2_79: begin
          r136_transform_384_545 <= insn_o_2_296_0;
          st_2 <= `S_2_488;
        end
        `S_2_488: begin
          r139_transform_385_546 <= insn_o_2_686_0;
          st_2 <= `S_2_492;
        end
        `S_2_492: begin
          sram_addr_2 <= 32'd4;
          sram_wdata_2 <= r139_transform_385_546;
          st_2 <= `S_2_496;
        end
        `S_2_496: begin
          sram_addr_2 <= 32'd5;
          st_2 <= `S_2_80;
        end
        `S_2_80: begin
          r144_transform_386_547 <= insn_o_2_305_0;
          st_2 <= `S_2_497;
        end
        `S_2_497: begin
          r147_transform_387_548 <= insn_o_2_698_0;
          st_2 <= `S_2_501;
        end
        `S_2_501: begin
          sram_addr_2 <= 32'd5;
          sram_wdata_2 <= r147_transform_387_548;
          st_2 <= `S_2_505;
        end
        `S_2_505: begin
          sram_addr_2 <= 32'd6;
          st_2 <= `S_2_82;
        end
        `S_2_82: begin
          r152_transform_388_549 <= insn_o_2_310_0;
          st_2 <= `S_2_506;
        end
        `S_2_506: begin
          r155_transform_389_550 <= insn_o_2_710_0;
          st_2 <= `S_2_510;
        end
        `S_2_510: begin
          sram_addr_2 <= 32'd6;
          sram_wdata_2 <= r155_transform_389_550;
          st_2 <= `S_2_514;
        end
        `S_2_514: begin
          sram_addr_2 <= 32'd7;
          st_2 <= `S_2_83;
        end
        `S_2_83: begin
          r160_transform_390_551 <= insn_o_2_318_0;
          st_2 <= `S_2_515;
        end
        `S_2_515: begin
          r163_transform_391_552 <= insn_o_2_722_0;
          st_2 <= `S_2_519;
        end
        `S_2_519: begin
          sram_addr_2 <= 32'd7;
          sram_wdata_2 <= r163_transform_391_552;
          st_2 <= `S_2_19;
        end
        `S_2_525: begin
          arg_177_561 <= x_224_554;
          st_2 <= `S_2_542;
        end
        `S_2_526: begin
          r4_s1_226_555 <= r1_ror32_17_178_565;
          st_2 <= `S_2_528;
        end
        `S_2_528: begin
          arg_187_566 <= x_224_554;
          st_2 <= `S_2_555;
        end
        `S_2_529: begin
          r6_s1_227_556 <= r1_ror32_19_188_570;
          st_2 <= `S_2_530;
        end
        `S_2_530: begin
          r3_s1_228_557 <= insn_o_2_745_0;
          st_2 <= `S_2_532;
        end
        `S_2_532: begin
          r8_s1_229_558 <= insn_o_2_748_0;
          st_2 <= `S_2_533;
        end
        `S_2_533: begin
          r2_s1_230_559 <= insn_o_2_750_0;
          st_2 <= `S_2_534;
        end
        `S_2_534: begin
          r1_s1_225_560 <= r2_s1_230_559;
          st_2 <= `S_2_369;
        end
        `S_2_542: begin
          r3_ror32_17_179_562 <= insn_o_2_761_0;
          st_2 <= `S_2_545;
        end
        `S_2_545: begin
          r6_ror32_17_180_563 <= insn_o_2_765_0;
          st_2 <= `S_2_546;
        end
        `S_2_546: begin
          r2_ror32_17_181_564 <= insn_o_2_767_0;
          st_2 <= `S_2_547;
        end
        `S_2_547: begin
          r1_ror32_17_178_565 <= r2_ror32_17_181_564;
          st_2 <= `S_2_526;
        end
        `S_2_555: begin
          r3_ror32_19_189_567 <= insn_o_2_778_0;
          st_2 <= `S_2_558;
        end
        `S_2_558: begin
          r6_ror32_19_190_568 <= insn_o_2_782_0;
          st_2 <= `S_2_559;
        end
        `S_2_559: begin
          r2_ror32_19_191_569 <= insn_o_2_784_0;
          st_2 <= `S_2_560;
        end
        `S_2_560: begin
          r1_ror32_19_188_570 <= r2_ror32_19_191_569;
          st_2 <= `S_2_529;
        end
        `S_2_567: begin
          arg_212_578 <= x_217_571;
          st_2 <= `S_2_584;
        end
        `S_2_568: begin
          r4_s0_219_572 <= r1_ror32_7_213_582;
          st_2 <= `S_2_570;
        end
        `S_2_570: begin
          arg_182_583 <= x_217_571;
          st_2 <= `S_2_597;
        end
        `S_2_571: begin
          r6_s0_220_573 <= r1_ror32_18_183_587;
          st_2 <= `S_2_572;
        end
        `S_2_572: begin
          r3_s0_221_574 <= insn_o_2_805_0;
          st_2 <= `S_2_574;
        end
        `S_2_574: begin
          r8_s0_222_575 <= insn_o_2_808_0;
          st_2 <= `S_2_575;
        end
        `S_2_575: begin
          r2_s0_223_576 <= insn_o_2_810_0;
          st_2 <= `S_2_576;
        end
        `S_2_576: begin
          r1_s0_218_577 <= r2_s0_223_576;
          st_2 <= `S_2_383;
        end
        `S_2_584: begin
          r3_ror32_7_214_579 <= insn_o_2_821_0;
          st_2 <= `S_2_587;
        end
        `S_2_587: begin
          r6_ror32_7_215_580 <= insn_o_2_825_0;
          st_2 <= `S_2_588;
        end
        `S_2_588: begin
          r2_ror32_7_216_581 <= insn_o_2_827_0;
          st_2 <= `S_2_589;
        end
        `S_2_589: begin
          r1_ror32_7_213_582 <= r2_ror32_7_216_581;
          st_2 <= `S_2_568;
        end
        `S_2_597: begin
          r3_ror32_18_184_584 <= insn_o_2_838_0;
          st_2 <= `S_2_600;
        end
        `S_2_600: begin
          r6_ror32_18_185_585 <= insn_o_2_842_0;
          st_2 <= `S_2_601;
        end
        `S_2_601: begin
          r2_ror32_18_186_586 <= insn_o_2_844_0;
          st_2 <= `S_2_602;
        end
        `S_2_602: begin
          r1_ror32_18_183_587 <= r2_ror32_18_186_586;
          st_2 <= `S_2_571;
        end
        `S_2_609: begin
          x_22_725 <= e_34_588;
          st_2 <= `S_2_882;
        end
        `S_2_610: begin
          r23_iterate_47_589 <= r1_e1_23_731;
          st_2 <= `S_2_611;
        end
        `S_2_611: begin
          r22_iterate_48_591 <= insn_o_2_859_0;
          st_2 <= `S_2_613;
        end
        `S_2_613: begin
          x_0_750 <= e_34_588;
          y_1_747 <= f_35_592;
          z_2_748 <= g_36_593;
          st_2 <= `S_2_937;
        end
        `S_2_614: begin
          r25_iterate_49_594 <= r3_Ch_3_753;
          st_2 <= `S_2_615;
        end
        `S_2_615: begin
          r21_iterate_50_595 <= insn_o_2_869_0;
          st_2 <= `S_2_618;
        end
        `S_2_618: begin
          sram_addr_222 <= idx_38_596;
          st_2 <= `S_2_86;
        end
        `S_2_86: begin
          r27_iterate_51_597 <= insn_o_2_327_0;
          st_2 <= `S_2_619;
        end
        `S_2_619: begin
          r20_iterate_52_598 <= insn_o_2_875_0;
          st_2 <= `S_2_622;
        end
        `S_2_622: begin
          sram_addr_223 <= idx_38_596;
          st_2 <= `S_2_87;
        end
        `S_2_87: begin
          r30_iterate_53_599 <= insn_o_2_330_0;
          st_2 <= `S_2_623;
        end
        `S_2_623: begin
          r19_iterate_54_600 <= insn_o_2_881_0;
          st_2 <= `S_2_624;
        end
        `S_2_624: begin
          r17_iterate_55_601 <= r19_iterate_54_600;
          st_2 <= `S_2_626;
        end
        `S_2_626: begin
          x_15_754 <= a_30_602;
          st_2 <= `S_2_947;
        end
        `S_2_627: begin
          r34_iterate_56_603 <= r1_e0_16_760;
          st_2 <= `S_2_629;
        end
        `S_2_629: begin
          x_7_776 <= a_30_602;
          y_8_777 <= b_31_604;
          z_9_780 <= c_32_605;
          st_2 <= `S_2_1002;
        end
        `S_2_630: begin
          r36_iterate_57_606 <= r3_Maj_10_783;
          st_2 <= `S_2_631;
        end
        `S_2_631: begin
          r33_iterate_58_607 <= insn_o_2_899_0;
          st_2 <= `S_2_632;
        end
        `S_2_632: begin
          r18_iterate_59_608 <= r33_iterate_58_607;
          st_2 <= `S_2_633;
        end
        `S_2_633: begin
          r38_iterate_60_610 <= insn_o_2_903_0;
          st_2 <= `S_2_634;
        end
        `S_2_634: begin
          d_33_609 <= r38_iterate_60_610;
          st_2 <= `S_2_635;
        end
        `S_2_635: begin
          r39_iterate_61_611 <= insn_o_2_907_0;
          st_2 <= `S_2_636;
        end
        `S_2_636: begin
          h_37_590 <= r39_iterate_61_611;
          st_2 <= `S_2_638;
        end
        `S_2_638: begin
          x_22_784 <= d_33_609;
          st_2 <= `S_2_1013;
        end
        `S_2_639: begin
          r44_iterate_62_612 <= r1_e1_23_790;
          st_2 <= `S_2_640;
        end
        `S_2_640: begin
          r43_iterate_63_613 <= insn_o_2_917_0;
          st_2 <= `S_2_642;
        end
        `S_2_642: begin
          x_0_809 <= d_33_609;
          y_1_806 <= e_34_588;
          z_2_807 <= f_35_592;
          st_2 <= `S_2_1068;
        end
        `S_2_643: begin
          r46_iterate_64_614 <= r3_Ch_3_812;
          st_2 <= `S_2_644;
        end
        `S_2_644: begin
          r42_iterate_65_615 <= insn_o_2_927_0;
          st_2 <= `S_2_646;
        end
        `S_2_646: begin
          r48_iterate_66_616 <= insn_o_2_930_0;
          st_2 <= `S_2_649;
        end
        `S_2_649: begin
          sram_addr_222 <= r48_iterate_66_616;
          st_2 <= `S_2_88;
        end
        `S_2_88: begin
          r50_iterate_67_617 <= insn_o_2_338_0;
          st_2 <= `S_2_650;
        end
        `S_2_650: begin
          r41_iterate_68_618 <= insn_o_2_936_0;
          st_2 <= `S_2_652;
        end
        `S_2_652: begin
          r53_iterate_69_619 <= insn_o_2_939_0;
          st_2 <= `S_2_655;
        end
        `S_2_655: begin
          sram_addr_223 <= r53_iterate_69_619;
          st_2 <= `S_2_90;
        end
        `S_2_90: begin
          r55_iterate_70_620 <= insn_o_2_341_0;
          st_2 <= `S_2_656;
        end
        `S_2_656: begin
          r40_iterate_71_621 <= insn_o_2_945_0;
          st_2 <= `S_2_657;
        end
        `S_2_657: begin
          r17_iterate_55_601 <= r40_iterate_71_621;
          st_2 <= `S_2_659;
        end
        `S_2_659: begin
          x_15_813 <= h_37_590;
          st_2 <= `S_2_1078;
        end
        `S_2_660: begin
          r59_iterate_72_622 <= r1_e0_16_819;
          st_2 <= `S_2_662;
        end
        `S_2_662: begin
          x_7_835 <= h_37_590;
          y_8_836 <= a_30_602;
          z_9_839 <= b_31_604;
          st_2 <= `S_2_1133;
        end
        `S_2_663: begin
          r61_iterate_73_623 <= r3_Maj_10_842;
          st_2 <= `S_2_664;
        end
        `S_2_664: begin
          r58_iterate_74_624 <= insn_o_2_963_0;
          st_2 <= `S_2_665;
        end
        `S_2_665: begin
          r18_iterate_59_608 <= r58_iterate_74_624;
          st_2 <= `S_2_666;
        end
        `S_2_666: begin
          r63_iterate_75_625 <= insn_o_2_967_0;
          st_2 <= `S_2_667;
        end
        `S_2_667: begin
          c_32_605 <= r63_iterate_75_625;
          st_2 <= `S_2_668;
        end
        `S_2_668: begin
          r64_iterate_76_626 <= insn_o_2_971_0;
          st_2 <= `S_2_669;
        end
        `S_2_669: begin
          g_36_593 <= r64_iterate_76_626;
          st_2 <= `S_2_671;
        end
        `S_2_671: begin
          x_22_843 <= c_32_605;
          st_2 <= `S_2_1144;
        end
        `S_2_672: begin
          r69_iterate_77_627 <= r1_e1_23_849;
          st_2 <= `S_2_673;
        end
        `S_2_673: begin
          r68_iterate_78_628 <= insn_o_2_981_0;
          st_2 <= `S_2_675;
        end
        `S_2_675: begin
          x_0_868 <= c_32_605;
          y_1_865 <= d_33_609;
          z_2_866 <= e_34_588;
          st_2 <= `S_2_1199;
        end
        `S_2_676: begin
          r71_iterate_79_629 <= r3_Ch_3_871;
          st_2 <= `S_2_677;
        end
        `S_2_677: begin
          r67_iterate_80_630 <= insn_o_2_991_0;
          st_2 <= `S_2_679;
        end
        `S_2_679: begin
          r73_iterate_81_631 <= insn_o_2_994_0;
          st_2 <= `S_2_682;
        end
        `S_2_682: begin
          sram_addr_222 <= r73_iterate_81_631;
          st_2 <= `S_2_91;
        end
        `S_2_91: begin
          r75_iterate_82_632 <= insn_o_2_349_0;
          st_2 <= `S_2_683;
        end
        `S_2_683: begin
          r66_iterate_83_633 <= insn_o_2_1000_0;
          st_2 <= `S_2_685;
        end
        `S_2_685: begin
          r78_iterate_84_634 <= insn_o_2_1003_0;
          st_2 <= `S_2_688;
        end
        `S_2_688: begin
          sram_addr_223 <= r78_iterate_84_634;
          st_2 <= `S_2_94;
        end
        `S_2_94: begin
          r80_iterate_85_635 <= insn_o_2_352_0;
          st_2 <= `S_2_689;
        end
        `S_2_689: begin
          r65_iterate_86_636 <= insn_o_2_1009_0;
          st_2 <= `S_2_690;
        end
        `S_2_690: begin
          r17_iterate_55_601 <= r65_iterate_86_636;
          st_2 <= `S_2_692;
        end
        `S_2_692: begin
          x_15_872 <= g_36_593;
          st_2 <= `S_2_1209;
        end
        `S_2_693: begin
          r84_iterate_87_637 <= r1_e0_16_878;
          st_2 <= `S_2_695;
        end
        `S_2_695: begin
          x_7_894 <= g_36_593;
          y_8_895 <= h_37_590;
          z_9_898 <= a_30_602;
          st_2 <= `S_2_1264;
        end
        `S_2_696: begin
          r86_iterate_88_638 <= r3_Maj_10_901;
          st_2 <= `S_2_697;
        end
        `S_2_697: begin
          r83_iterate_89_639 <= insn_o_2_1027_0;
          st_2 <= `S_2_698;
        end
        `S_2_698: begin
          r18_iterate_59_608 <= r83_iterate_89_639;
          st_2 <= `S_2_699;
        end
        `S_2_699: begin
          r88_iterate_90_640 <= insn_o_2_1031_0;
          st_2 <= `S_2_700;
        end
        `S_2_700: begin
          b_31_604 <= r88_iterate_90_640;
          st_2 <= `S_2_701;
        end
        `S_2_701: begin
          r89_iterate_91_641 <= insn_o_2_1035_0;
          st_2 <= `S_2_702;
        end
        `S_2_702: begin
          f_35_592 <= r89_iterate_91_641;
          st_2 <= `S_2_704;
        end
        `S_2_704: begin
          x_22_902 <= b_31_604;
          st_2 <= `S_2_1275;
        end
        `S_2_705: begin
          r94_iterate_92_642 <= r1_e1_23_908;
          st_2 <= `S_2_706;
        end
        `S_2_706: begin
          r93_iterate_93_643 <= insn_o_2_1045_0;
          st_2 <= `S_2_708;
        end
        `S_2_708: begin
          x_0_927 <= b_31_604;
          y_1_924 <= c_32_605;
          z_2_925 <= d_33_609;
          st_2 <= `S_2_1330;
        end
        `S_2_709: begin
          r96_iterate_94_644 <= r3_Ch_3_930;
          st_2 <= `S_2_710;
        end
        `S_2_710: begin
          r92_iterate_95_645 <= insn_o_2_1055_0;
          st_2 <= `S_2_712;
        end
        `S_2_712: begin
          r98_iterate_96_646 <= insn_o_2_1058_0;
          st_2 <= `S_2_715;
        end
        `S_2_715: begin
          sram_addr_222 <= r98_iterate_96_646;
          st_2 <= `S_2_95;
        end
        `S_2_95: begin
          r100_iterate_97_647 <= insn_o_2_360_0;
          st_2 <= `S_2_716;
        end
        `S_2_716: begin
          r91_iterate_98_648 <= insn_o_2_1064_0;
          st_2 <= `S_2_718;
        end
        `S_2_718: begin
          r103_iterate_99_649 <= insn_o_2_1067_0;
          st_2 <= `S_2_721;
        end
        `S_2_721: begin
          sram_addr_223 <= r103_iterate_99_649;
          st_2 <= `S_2_96;
        end
        `S_2_96: begin
          r105_iterate_100_650 <= insn_o_2_363_0;
          st_2 <= `S_2_722;
        end
        `S_2_722: begin
          r90_iterate_101_651 <= insn_o_2_1073_0;
          st_2 <= `S_2_723;
        end
        `S_2_723: begin
          r17_iterate_55_601 <= r90_iterate_101_651;
          st_2 <= `S_2_725;
        end
        `S_2_725: begin
          x_15_931 <= f_35_592;
          st_2 <= `S_2_1340;
        end
        `S_2_726: begin
          r109_iterate_102_652 <= r1_e0_16_937;
          st_2 <= `S_2_728;
        end
        `S_2_728: begin
          x_7_953 <= f_35_592;
          y_8_954 <= g_36_593;
          z_9_957 <= h_37_590;
          st_2 <= `S_2_1395;
        end
        `S_2_729: begin
          r111_iterate_103_653 <= r3_Maj_10_960;
          st_2 <= `S_2_730;
        end
        `S_2_730: begin
          r108_iterate_104_654 <= insn_o_2_1091_0;
          st_2 <= `S_2_731;
        end
        `S_2_731: begin
          r18_iterate_59_608 <= r108_iterate_104_654;
          st_2 <= `S_2_732;
        end
        `S_2_732: begin
          r113_iterate_105_655 <= insn_o_2_1095_0;
          st_2 <= `S_2_733;
        end
        `S_2_733: begin
          a_30_602 <= r113_iterate_105_655;
          st_2 <= `S_2_734;
        end
        `S_2_734: begin
          r114_iterate_106_656 <= insn_o_2_1099_0;
          st_2 <= `S_2_735;
        end
        `S_2_735: begin
          e_34_588 <= r114_iterate_106_656;
          st_2 <= `S_2_737;
        end
        `S_2_737: begin
          x_22_961 <= a_30_602;
          st_2 <= `S_2_1406;
        end
        `S_2_738: begin
          r119_iterate_107_657 <= r1_e1_23_967;
          st_2 <= `S_2_739;
        end
        `S_2_739: begin
          r118_iterate_108_658 <= insn_o_2_1109_0;
          st_2 <= `S_2_741;
        end
        `S_2_741: begin
          x_0_986 <= a_30_602;
          y_1_983 <= b_31_604;
          z_2_984 <= c_32_605;
          st_2 <= `S_2_1461;
        end
        `S_2_742: begin
          r121_iterate_109_659 <= r3_Ch_3_989;
          st_2 <= `S_2_743;
        end
        `S_2_743: begin
          r117_iterate_110_660 <= insn_o_2_1119_0;
          st_2 <= `S_2_745;
        end
        `S_2_745: begin
          r123_iterate_111_661 <= insn_o_2_1122_0;
          st_2 <= `S_2_748;
        end
        `S_2_748: begin
          sram_addr_222 <= r123_iterate_111_661;
          st_2 <= `S_2_98;
        end
        `S_2_98: begin
          r125_iterate_112_662 <= insn_o_2_371_0;
          st_2 <= `S_2_749;
        end
        `S_2_749: begin
          r116_iterate_113_663 <= insn_o_2_1128_0;
          st_2 <= `S_2_751;
        end
        `S_2_751: begin
          r128_iterate_114_664 <= insn_o_2_1131_0;
          st_2 <= `S_2_754;
        end
        `S_2_754: begin
          sram_addr_223 <= r128_iterate_114_664;
          st_2 <= `S_2_99;
        end
        `S_2_99: begin
          r130_iterate_115_665 <= insn_o_2_374_0;
          st_2 <= `S_2_755;
        end
        `S_2_755: begin
          r115_iterate_116_666 <= insn_o_2_1137_0;
          st_2 <= `S_2_756;
        end
        `S_2_756: begin
          r17_iterate_55_601 <= r115_iterate_116_666;
          st_2 <= `S_2_758;
        end
        `S_2_758: begin
          x_15_990 <= e_34_588;
          st_2 <= `S_2_1471;
        end
        `S_2_759: begin
          r134_iterate_117_667 <= r1_e0_16_996;
          st_2 <= `S_2_761;
        end
        `S_2_761: begin
          x_7_1012 <= e_34_588;
          y_8_1013 <= f_35_592;
          z_9_1016 <= g_36_593;
          st_2 <= `S_2_1526;
        end
        `S_2_762: begin
          r136_iterate_118_668 <= r3_Maj_10_1019;
          st_2 <= `S_2_763;
        end
        `S_2_763: begin
          r133_iterate_119_669 <= insn_o_2_1155_0;
          st_2 <= `S_2_764;
        end
        `S_2_764: begin
          r18_iterate_59_608 <= r133_iterate_119_669;
          st_2 <= `S_2_765;
        end
        `S_2_765: begin
          r138_iterate_120_670 <= insn_o_2_1159_0;
          st_2 <= `S_2_766;
        end
        `S_2_766: begin
          h_37_590 <= r138_iterate_120_670;
          st_2 <= `S_2_767;
        end
        `S_2_767: begin
          r139_iterate_121_671 <= insn_o_2_1163_0;
          st_2 <= `S_2_768;
        end
        `S_2_768: begin
          d_33_609 <= r139_iterate_121_671;
          st_2 <= `S_2_770;
        end
        `S_2_770: begin
          x_22_1020 <= h_37_590;
          st_2 <= `S_2_1537;
        end
        `S_2_771: begin
          r144_iterate_122_672 <= r1_e1_23_1026;
          st_2 <= `S_2_772;
        end
        `S_2_772: begin
          r143_iterate_123_673 <= insn_o_2_1173_0;
          st_2 <= `S_2_774;
        end
        `S_2_774: begin
          x_0_1045 <= h_37_590;
          y_1_1042 <= a_30_602;
          z_2_1043 <= b_31_604;
          st_2 <= `S_2_1592;
        end
        `S_2_775: begin
          r146_iterate_124_674 <= r3_Ch_3_1048;
          st_2 <= `S_2_776;
        end
        `S_2_776: begin
          r142_iterate_125_675 <= insn_o_2_1183_0;
          st_2 <= `S_2_778;
        end
        `S_2_778: begin
          r148_iterate_126_676 <= insn_o_2_1186_0;
          st_2 <= `S_2_781;
        end
        `S_2_781: begin
          sram_addr_222 <= r148_iterate_126_676;
          st_2 <= `S_2_102;
        end
        `S_2_102: begin
          r150_iterate_127_677 <= insn_o_2_384_0;
          st_2 <= `S_2_782;
        end
        `S_2_782: begin
          r141_iterate_128_678 <= insn_o_2_1192_0;
          st_2 <= `S_2_784;
        end
        `S_2_784: begin
          r153_iterate_129_679 <= insn_o_2_1195_0;
          st_2 <= `S_2_787;
        end
        `S_2_787: begin
          sram_addr_223 <= r153_iterate_129_679;
          st_2 <= `S_2_103;
        end
        `S_2_103: begin
          r155_iterate_130_680 <= insn_o_2_388_0;
          st_2 <= `S_2_788;
        end
        `S_2_788: begin
          r140_iterate_131_681 <= insn_o_2_1201_0;
          st_2 <= `S_2_789;
        end
        `S_2_789: begin
          r17_iterate_55_601 <= r140_iterate_131_681;
          st_2 <= `S_2_791;
        end
        `S_2_791: begin
          x_15_1049 <= d_33_609;
          st_2 <= `S_2_1602;
        end
        `S_2_792: begin
          r159_iterate_132_682 <= r1_e0_16_1055;
          st_2 <= `S_2_794;
        end
        `S_2_794: begin
          x_7_1071 <= d_33_609;
          y_8_1072 <= e_34_588;
          z_9_1075 <= f_35_592;
          st_2 <= `S_2_1657;
        end
        `S_2_795: begin
          r161_iterate_133_683 <= r3_Maj_10_1078;
          st_2 <= `S_2_796;
        end
        `S_2_796: begin
          r158_iterate_134_684 <= insn_o_2_1219_0;
          st_2 <= `S_2_797;
        end
        `S_2_797: begin
          r18_iterate_59_608 <= r158_iterate_134_684;
          st_2 <= `S_2_798;
        end
        `S_2_798: begin
          r163_iterate_135_685 <= insn_o_2_1223_0;
          st_2 <= `S_2_799;
        end
        `S_2_799: begin
          g_36_593 <= r163_iterate_135_685;
          st_2 <= `S_2_800;
        end
        `S_2_800: begin
          r164_iterate_136_686 <= insn_o_2_1227_0;
          st_2 <= `S_2_801;
        end
        `S_2_801: begin
          c_32_605 <= r164_iterate_136_686;
          st_2 <= `S_2_803;
        end
        `S_2_803: begin
          x_22_1079 <= g_36_593;
          st_2 <= `S_2_1668;
        end
        `S_2_804: begin
          r169_iterate_137_687 <= r1_e1_23_1085;
          st_2 <= `S_2_805;
        end
        `S_2_805: begin
          r168_iterate_138_688 <= insn_o_2_1237_0;
          st_2 <= `S_2_807;
        end
        `S_2_807: begin
          x_0_1104 <= g_36_593;
          y_1_1101 <= h_37_590;
          z_2_1102 <= a_30_602;
          st_2 <= `S_2_1723;
        end
        `S_2_808: begin
          r171_iterate_139_689 <= r3_Ch_3_1107;
          st_2 <= `S_2_809;
        end
        `S_2_809: begin
          r167_iterate_140_690 <= insn_o_2_1247_0;
          st_2 <= `S_2_811;
        end
        `S_2_811: begin
          r173_iterate_141_691 <= insn_o_2_1250_0;
          st_2 <= `S_2_814;
        end
        `S_2_814: begin
          sram_addr_222 <= r173_iterate_141_691;
          st_2 <= `S_2_104;
        end
        `S_2_104: begin
          r175_iterate_142_692 <= insn_o_2_391_0;
          st_2 <= `S_2_815;
        end
        `S_2_815: begin
          r166_iterate_143_693 <= insn_o_2_1256_0;
          st_2 <= `S_2_817;
        end
        `S_2_817: begin
          r178_iterate_144_694 <= insn_o_2_1259_0;
          st_2 <= `S_2_820;
        end
        `S_2_820: begin
          sram_addr_223 <= r178_iterate_144_694;
          st_2 <= `S_2_106;
        end
        `S_2_106: begin
          r180_iterate_145_695 <= insn_o_2_395_0;
          st_2 <= `S_2_821;
        end
        `S_2_821: begin
          r165_iterate_146_696 <= insn_o_2_1265_0;
          st_2 <= `S_2_822;
        end
        `S_2_822: begin
          r17_iterate_55_601 <= r165_iterate_146_696;
          st_2 <= `S_2_824;
        end
        `S_2_824: begin
          x_15_1108 <= c_32_605;
          st_2 <= `S_2_1733;
        end
        `S_2_825: begin
          r184_iterate_147_697 <= r1_e0_16_1114;
          st_2 <= `S_2_827;
        end
        `S_2_827: begin
          x_7_1130 <= c_32_605;
          y_8_1131 <= d_33_609;
          z_9_1134 <= e_34_588;
          st_2 <= `S_2_1788;
        end
        `S_2_828: begin
          r186_iterate_148_698 <= r3_Maj_10_1137;
          st_2 <= `S_2_829;
        end
        `S_2_829: begin
          r183_iterate_149_699 <= insn_o_2_1283_0;
          st_2 <= `S_2_830;
        end
        `S_2_830: begin
          r18_iterate_59_608 <= r183_iterate_149_699;
          st_2 <= `S_2_831;
        end
        `S_2_831: begin
          r188_iterate_150_700 <= insn_o_2_1287_0;
          st_2 <= `S_2_832;
        end
        `S_2_832: begin
          f_35_592 <= r188_iterate_150_700;
          st_2 <= `S_2_833;
        end
        `S_2_833: begin
          r189_iterate_151_701 <= insn_o_2_1291_0;
          st_2 <= `S_2_834;
        end
        `S_2_834: begin
          b_31_604 <= r189_iterate_151_701;
          st_2 <= `S_2_836;
        end
        `S_2_836: begin
          x_22_1138 <= f_35_592;
          st_2 <= `S_2_1799;
        end
        `S_2_837: begin
          r194_iterate_152_702 <= r1_e1_23_1144;
          st_2 <= `S_2_838;
        end
        `S_2_838: begin
          r193_iterate_153_703 <= insn_o_2_1301_0;
          st_2 <= `S_2_840;
        end
        `S_2_840: begin
          x_0_1163 <= f_35_592;
          y_1_1160 <= g_36_593;
          z_2_1161 <= h_37_590;
          st_2 <= `S_2_1854;
        end
        `S_2_841: begin
          r196_iterate_154_704 <= r3_Ch_3_1166;
          st_2 <= `S_2_842;
        end
        `S_2_842: begin
          r192_iterate_155_705 <= insn_o_2_1311_0;
          st_2 <= `S_2_844;
        end
        `S_2_844: begin
          r198_iterate_156_706 <= insn_o_2_1314_0;
          st_2 <= `S_2_847;
        end
        `S_2_847: begin
          sram_addr_222 <= r198_iterate_156_706;
          st_2 <= `S_2_107;
        end
        `S_2_107: begin
          r200_iterate_157_707 <= insn_o_2_398_0;
          st_2 <= `S_2_848;
        end
        `S_2_848: begin
          r191_iterate_158_708 <= insn_o_2_1320_0;
          st_2 <= `S_2_850;
        end
        `S_2_850: begin
          r203_iterate_159_709 <= insn_o_2_1323_0;
          st_2 <= `S_2_853;
        end
        `S_2_853: begin
          sram_addr_223 <= r203_iterate_159_709;
          st_2 <= `S_2_110;
        end
        `S_2_110: begin
          r205_iterate_160_710 <= insn_o_2_402_0;
          st_2 <= `S_2_854;
        end
        `S_2_854: begin
          r190_iterate_161_711 <= insn_o_2_1329_0;
          st_2 <= `S_2_855;
        end
        `S_2_855: begin
          r17_iterate_55_601 <= r190_iterate_161_711;
          st_2 <= `S_2_857;
        end
        `S_2_857: begin
          x_15_1167 <= b_31_604;
          st_2 <= `S_2_1864;
        end
        `S_2_858: begin
          r209_iterate_162_712 <= r1_e0_16_1173;
          st_2 <= `S_2_860;
        end
        `S_2_860: begin
          x_7_1189 <= b_31_604;
          y_8_1190 <= c_32_605;
          z_9_1193 <= d_33_609;
          st_2 <= `S_2_1919;
        end
        `S_2_861: begin
          r211_iterate_163_713 <= r3_Maj_10_1196;
          st_2 <= `S_2_862;
        end
        `S_2_862: begin
          r208_iterate_164_714 <= insn_o_2_1347_0;
          st_2 <= `S_2_863;
        end
        `S_2_863: begin
          r18_iterate_59_608 <= r208_iterate_164_714;
          st_2 <= `S_2_864;
        end
        `S_2_864: begin
          r213_iterate_165_715 <= insn_o_2_1351_0;
          st_2 <= `S_2_865;
        end
        `S_2_865: begin
          e_34_588 <= r213_iterate_165_715;
          st_2 <= `S_2_866;
        end
        `S_2_866: begin
          r214_iterate_166_716 <= insn_o_2_1355_0;
          st_2 <= `S_2_867;
        end
        `S_2_867: begin
          a_30_602 <= r214_iterate_166_716;
          st_2 <= `S_2_868;
        end
        `S_2_868: begin
          r9_iterate_39_717 <= a_30_602;
          st_2 <= `S_2_869;
        end
        `S_2_869: begin
          r10_iterate_40_718 <= b_31_604;
          st_2 <= `S_2_870;
        end
        `S_2_870: begin
          r11_iterate_41_719 <= c_32_605;
          st_2 <= `S_2_871;
        end
        `S_2_871: begin
          r12_iterate_42_720 <= d_33_609;
          st_2 <= `S_2_872;
        end
        `S_2_872: begin
          r13_iterate_43_721 <= e_34_588;
          st_2 <= `S_2_873;
        end
        `S_2_873: begin
          r14_iterate_44_722 <= f_35_592;
          st_2 <= `S_2_874;
        end
        `S_2_874: begin
          r15_iterate_45_723 <= g_36_593;
          st_2 <= `S_2_875;
        end
        `S_2_875: begin
          r16_iterate_46_724 <= h_37_590;
          st_2 <= `S_2_443;
        end
        `S_2_882: begin
          arg_207_732 <= x_22_725;
          st_2 <= `S_2_900;
        end
        `S_2_883: begin
          r4_e1_24_726 <= r1_ror32_6_208_736;
          st_2 <= `S_2_885;
        end
        `S_2_885: begin
          arg_167_737 <= x_22_725;
          st_2 <= `S_2_913;
        end
        `S_2_886: begin
          r6_e1_25_727 <= r1_ror32_11_168_741;
          st_2 <= `S_2_887;
        end
        `S_2_887: begin
          r3_e1_26_728 <= insn_o_2_1392_0;
          st_2 <= `S_2_889;
        end
        `S_2_889: begin
          arg_202_742 <= x_22_725;
          st_2 <= `S_2_926;
        end
        `S_2_890: begin
          r8_e1_27_729 <= r1_ror32_25_203_746;
          st_2 <= `S_2_891;
        end
        `S_2_891: begin
          r2_e1_28_730 <= insn_o_2_1400_0;
          st_2 <= `S_2_892;
        end
        `S_2_892: begin
          r1_e1_23_731 <= r2_e1_28_730;
          st_2 <= `S_2_610;
        end
        `S_2_900: begin
          r3_ror32_6_209_733 <= insn_o_2_1411_0;
          st_2 <= `S_2_903;
        end
        `S_2_903: begin
          r6_ror32_6_210_734 <= insn_o_2_1415_0;
          st_2 <= `S_2_904;
        end
        `S_2_904: begin
          r2_ror32_6_211_735 <= insn_o_2_1417_0;
          st_2 <= `S_2_905;
        end
        `S_2_905: begin
          r1_ror32_6_208_736 <= r2_ror32_6_211_735;
          st_2 <= `S_2_883;
        end
        `S_2_913: begin
          r3_ror32_11_169_738 <= insn_o_2_1428_0;
          st_2 <= `S_2_916;
        end
        `S_2_916: begin
          r6_ror32_11_170_739 <= insn_o_2_1432_0;
          st_2 <= `S_2_917;
        end
        `S_2_917: begin
          r2_ror32_11_171_740 <= insn_o_2_1434_0;
          st_2 <= `S_2_918;
        end
        `S_2_918: begin
          r1_ror32_11_168_741 <= r2_ror32_11_171_740;
          st_2 <= `S_2_886;
        end
        `S_2_926: begin
          r3_ror32_25_204_743 <= insn_o_2_1445_0;
          st_2 <= `S_2_929;
        end
        `S_2_929: begin
          r6_ror32_25_205_744 <= insn_o_2_1449_0;
          st_2 <= `S_2_930;
        end
        `S_2_930: begin
          r2_ror32_25_206_745 <= insn_o_2_1451_0;
          st_2 <= `S_2_931;
        end
        `S_2_931: begin
          r1_ror32_25_203_746 <= r2_ror32_25_206_745;
          st_2 <= `S_2_890;
        end
        `S_2_937: begin
          r6_Ch_4_749 <= insn_o_2_1460_0;
          st_2 <= `S_2_938;
        end
        `S_2_938: begin
          r5_Ch_5_751 <= insn_o_2_1462_0;
          st_2 <= `S_2_939;
        end
        `S_2_939: begin
          r4_Ch_6_752 <= insn_o_2_1464_0;
          st_2 <= `S_2_940;
        end
        `S_2_940: begin
          r3_Ch_3_753 <= r4_Ch_6_752;
          st_2 <= `S_2_614;
        end
        `S_2_947: begin
          arg_192_761 <= x_15_754;
          st_2 <= `S_2_965;
        end
        `S_2_948: begin
          r4_e0_17_755 <= r1_ror32_2_193_765;
          st_2 <= `S_2_950;
        end
        `S_2_950: begin
          arg_172_766 <= x_15_754;
          st_2 <= `S_2_978;
        end
        `S_2_951: begin
          r6_e0_18_756 <= r1_ror32_13_173_770;
          st_2 <= `S_2_952;
        end
        `S_2_952: begin
          r3_e0_19_757 <= insn_o_2_1485_0;
          st_2 <= `S_2_954;
        end
        `S_2_954: begin
          arg_197_771 <= x_15_754;
          st_2 <= `S_2_991;
        end
        `S_2_955: begin
          r8_e0_20_758 <= r1_ror32_22_198_775;
          st_2 <= `S_2_956;
        end
        `S_2_956: begin
          r2_e0_21_759 <= insn_o_2_1493_0;
          st_2 <= `S_2_957;
        end
        `S_2_957: begin
          r1_e0_16_760 <= r2_e0_21_759;
          st_2 <= `S_2_627;
        end
        `S_2_965: begin
          r3_ror32_2_194_762 <= insn_o_2_1504_0;
          st_2 <= `S_2_968;
        end
        `S_2_968: begin
          r6_ror32_2_195_763 <= insn_o_2_1508_0;
          st_2 <= `S_2_969;
        end
        `S_2_969: begin
          r2_ror32_2_196_764 <= insn_o_2_1510_0;
          st_2 <= `S_2_970;
        end
        `S_2_970: begin
          r1_ror32_2_193_765 <= r2_ror32_2_196_764;
          st_2 <= `S_2_948;
        end
        `S_2_978: begin
          r3_ror32_13_174_767 <= insn_o_2_1521_0;
          st_2 <= `S_2_981;
        end
        `S_2_981: begin
          r6_ror32_13_175_768 <= insn_o_2_1525_0;
          st_2 <= `S_2_982;
        end
        `S_2_982: begin
          r2_ror32_13_176_769 <= insn_o_2_1527_0;
          st_2 <= `S_2_983;
        end
        `S_2_983: begin
          r1_ror32_13_173_770 <= r2_ror32_13_176_769;
          st_2 <= `S_2_951;
        end
        `S_2_991: begin
          r3_ror32_22_199_772 <= insn_o_2_1538_0;
          st_2 <= `S_2_994;
        end
        `S_2_994: begin
          r6_ror32_22_200_773 <= insn_o_2_1542_0;
          st_2 <= `S_2_995;
        end
        `S_2_995: begin
          r2_ror32_22_201_774 <= insn_o_2_1544_0;
          st_2 <= `S_2_996;
        end
        `S_2_996: begin
          r1_ror32_22_198_775 <= r2_ror32_22_201_774;
          st_2 <= `S_2_955;
        end
        `S_2_1002: begin
          r5_Maj_11_778 <= insn_o_2_1553_0;
          st_2 <= `S_2_1003;
        end
        `S_2_1003: begin
          r7_Maj_12_779 <= insn_o_2_1555_0;
          st_2 <= `S_2_1004;
        end
        `S_2_1004: begin
          r6_Maj_13_781 <= insn_o_2_1557_0;
          st_2 <= `S_2_1005;
        end
        `S_2_1005: begin
          r4_Maj_14_782 <= insn_o_2_1559_0;
          st_2 <= `S_2_1006;
        end
        `S_2_1006: begin
          r3_Maj_10_783 <= r4_Maj_14_782;
          st_2 <= `S_2_630;
        end
        `S_2_1013: begin
          arg_207_791 <= x_22_784;
          st_2 <= `S_2_1031;
        end
        `S_2_1014: begin
          r4_e1_24_785 <= r1_ror32_6_208_795;
          st_2 <= `S_2_1016;
        end
        `S_2_1016: begin
          arg_167_796 <= x_22_784;
          st_2 <= `S_2_1044;
        end
        `S_2_1017: begin
          r6_e1_25_786 <= r1_ror32_11_168_800;
          st_2 <= `S_2_1018;
        end
        `S_2_1018: begin
          r3_e1_26_787 <= insn_o_2_1580_0;
          st_2 <= `S_2_1020;
        end
        `S_2_1020: begin
          arg_202_801 <= x_22_784;
          st_2 <= `S_2_1057;
        end
        `S_2_1021: begin
          r8_e1_27_788 <= r1_ror32_25_203_805;
          st_2 <= `S_2_1022;
        end
        `S_2_1022: begin
          r2_e1_28_789 <= insn_o_2_1588_0;
          st_2 <= `S_2_1023;
        end
        `S_2_1023: begin
          r1_e1_23_790 <= r2_e1_28_789;
          st_2 <= `S_2_639;
        end
        `S_2_1031: begin
          r3_ror32_6_209_792 <= insn_o_2_1599_0;
          st_2 <= `S_2_1034;
        end
        `S_2_1034: begin
          r6_ror32_6_210_793 <= insn_o_2_1603_0;
          st_2 <= `S_2_1035;
        end
        `S_2_1035: begin
          r2_ror32_6_211_794 <= insn_o_2_1605_0;
          st_2 <= `S_2_1036;
        end
        `S_2_1036: begin
          r1_ror32_6_208_795 <= r2_ror32_6_211_794;
          st_2 <= `S_2_1014;
        end
        `S_2_1044: begin
          r3_ror32_11_169_797 <= insn_o_2_1616_0;
          st_2 <= `S_2_1047;
        end
        `S_2_1047: begin
          r6_ror32_11_170_798 <= insn_o_2_1620_0;
          st_2 <= `S_2_1048;
        end
        `S_2_1048: begin
          r2_ror32_11_171_799 <= insn_o_2_1622_0;
          st_2 <= `S_2_1049;
        end
        `S_2_1049: begin
          r1_ror32_11_168_800 <= r2_ror32_11_171_799;
          st_2 <= `S_2_1017;
        end
        `S_2_1057: begin
          r3_ror32_25_204_802 <= insn_o_2_1633_0;
          st_2 <= `S_2_1060;
        end
        `S_2_1060: begin
          r6_ror32_25_205_803 <= insn_o_2_1637_0;
          st_2 <= `S_2_1061;
        end
        `S_2_1061: begin
          r2_ror32_25_206_804 <= insn_o_2_1639_0;
          st_2 <= `S_2_1062;
        end
        `S_2_1062: begin
          r1_ror32_25_203_805 <= r2_ror32_25_206_804;
          st_2 <= `S_2_1021;
        end
        `S_2_1068: begin
          r6_Ch_4_808 <= insn_o_2_1648_0;
          st_2 <= `S_2_1069;
        end
        `S_2_1069: begin
          r5_Ch_5_810 <= insn_o_2_1650_0;
          st_2 <= `S_2_1070;
        end
        `S_2_1070: begin
          r4_Ch_6_811 <= insn_o_2_1652_0;
          st_2 <= `S_2_1071;
        end
        `S_2_1071: begin
          r3_Ch_3_812 <= r4_Ch_6_811;
          st_2 <= `S_2_643;
        end
        `S_2_1078: begin
          arg_192_820 <= x_15_813;
          st_2 <= `S_2_1096;
        end
        `S_2_1079: begin
          r4_e0_17_814 <= r1_ror32_2_193_824;
          st_2 <= `S_2_1081;
        end
        `S_2_1081: begin
          arg_172_825 <= x_15_813;
          st_2 <= `S_2_1109;
        end
        `S_2_1082: begin
          r6_e0_18_815 <= r1_ror32_13_173_829;
          st_2 <= `S_2_1083;
        end
        `S_2_1083: begin
          r3_e0_19_816 <= insn_o_2_1673_0;
          st_2 <= `S_2_1085;
        end
        `S_2_1085: begin
          arg_197_830 <= x_15_813;
          st_2 <= `S_2_1122;
        end
        `S_2_1086: begin
          r8_e0_20_817 <= r1_ror32_22_198_834;
          st_2 <= `S_2_1087;
        end
        `S_2_1087: begin
          r2_e0_21_818 <= insn_o_2_1681_0;
          st_2 <= `S_2_1088;
        end
        `S_2_1088: begin
          r1_e0_16_819 <= r2_e0_21_818;
          st_2 <= `S_2_660;
        end
        `S_2_1096: begin
          r3_ror32_2_194_821 <= insn_o_2_1692_0;
          st_2 <= `S_2_1099;
        end
        `S_2_1099: begin
          r6_ror32_2_195_822 <= insn_o_2_1696_0;
          st_2 <= `S_2_1100;
        end
        `S_2_1100: begin
          r2_ror32_2_196_823 <= insn_o_2_1698_0;
          st_2 <= `S_2_1101;
        end
        `S_2_1101: begin
          r1_ror32_2_193_824 <= r2_ror32_2_196_823;
          st_2 <= `S_2_1079;
        end
        `S_2_1109: begin
          r3_ror32_13_174_826 <= insn_o_2_1709_0;
          st_2 <= `S_2_1112;
        end
        `S_2_1112: begin
          r6_ror32_13_175_827 <= insn_o_2_1713_0;
          st_2 <= `S_2_1113;
        end
        `S_2_1113: begin
          r2_ror32_13_176_828 <= insn_o_2_1715_0;
          st_2 <= `S_2_1114;
        end
        `S_2_1114: begin
          r1_ror32_13_173_829 <= r2_ror32_13_176_828;
          st_2 <= `S_2_1082;
        end
        `S_2_1122: begin
          r3_ror32_22_199_831 <= insn_o_2_1726_0;
          st_2 <= `S_2_1125;
        end
        `S_2_1125: begin
          r6_ror32_22_200_832 <= insn_o_2_1730_0;
          st_2 <= `S_2_1126;
        end
        `S_2_1126: begin
          r2_ror32_22_201_833 <= insn_o_2_1732_0;
          st_2 <= `S_2_1127;
        end
        `S_2_1127: begin
          r1_ror32_22_198_834 <= r2_ror32_22_201_833;
          st_2 <= `S_2_1086;
        end
        `S_2_1133: begin
          r5_Maj_11_837 <= insn_o_2_1741_0;
          st_2 <= `S_2_1134;
        end
        `S_2_1134: begin
          r7_Maj_12_838 <= insn_o_2_1743_0;
          st_2 <= `S_2_1135;
        end
        `S_2_1135: begin
          r6_Maj_13_840 <= insn_o_2_1745_0;
          st_2 <= `S_2_1136;
        end
        `S_2_1136: begin
          r4_Maj_14_841 <= insn_o_2_1747_0;
          st_2 <= `S_2_1137;
        end
        `S_2_1137: begin
          r3_Maj_10_842 <= r4_Maj_14_841;
          st_2 <= `S_2_663;
        end
        `S_2_1144: begin
          arg_207_850 <= x_22_843;
          st_2 <= `S_2_1162;
        end
        `S_2_1145: begin
          r4_e1_24_844 <= r1_ror32_6_208_854;
          st_2 <= `S_2_1147;
        end
        `S_2_1147: begin
          arg_167_855 <= x_22_843;
          st_2 <= `S_2_1175;
        end
        `S_2_1148: begin
          r6_e1_25_845 <= r1_ror32_11_168_859;
          st_2 <= `S_2_1149;
        end
        `S_2_1149: begin
          r3_e1_26_846 <= insn_o_2_1768_0;
          st_2 <= `S_2_1151;
        end
        `S_2_1151: begin
          arg_202_860 <= x_22_843;
          st_2 <= `S_2_1188;
        end
        `S_2_1152: begin
          r8_e1_27_847 <= r1_ror32_25_203_864;
          st_2 <= `S_2_1153;
        end
        `S_2_1153: begin
          r2_e1_28_848 <= insn_o_2_1776_0;
          st_2 <= `S_2_1154;
        end
        `S_2_1154: begin
          r1_e1_23_849 <= r2_e1_28_848;
          st_2 <= `S_2_672;
        end
        `S_2_1162: begin
          r3_ror32_6_209_851 <= insn_o_2_1787_0;
          st_2 <= `S_2_1165;
        end
        `S_2_1165: begin
          r6_ror32_6_210_852 <= insn_o_2_1791_0;
          st_2 <= `S_2_1166;
        end
        `S_2_1166: begin
          r2_ror32_6_211_853 <= insn_o_2_1793_0;
          st_2 <= `S_2_1167;
        end
        `S_2_1167: begin
          r1_ror32_6_208_854 <= r2_ror32_6_211_853;
          st_2 <= `S_2_1145;
        end
        `S_2_1175: begin
          r3_ror32_11_169_856 <= insn_o_2_1804_0;
          st_2 <= `S_2_1178;
        end
        `S_2_1178: begin
          r6_ror32_11_170_857 <= insn_o_2_1808_0;
          st_2 <= `S_2_1179;
        end
        `S_2_1179: begin
          r2_ror32_11_171_858 <= insn_o_2_1810_0;
          st_2 <= `S_2_1180;
        end
        `S_2_1180: begin
          r1_ror32_11_168_859 <= r2_ror32_11_171_858;
          st_2 <= `S_2_1148;
        end
        `S_2_1188: begin
          r3_ror32_25_204_861 <= insn_o_2_1821_0;
          st_2 <= `S_2_1191;
        end
        `S_2_1191: begin
          r6_ror32_25_205_862 <= insn_o_2_1825_0;
          st_2 <= `S_2_1192;
        end
        `S_2_1192: begin
          r2_ror32_25_206_863 <= insn_o_2_1827_0;
          st_2 <= `S_2_1193;
        end
        `S_2_1193: begin
          r1_ror32_25_203_864 <= r2_ror32_25_206_863;
          st_2 <= `S_2_1152;
        end
        `S_2_1199: begin
          r6_Ch_4_867 <= insn_o_2_1836_0;
          st_2 <= `S_2_1200;
        end
        `S_2_1200: begin
          r5_Ch_5_869 <= insn_o_2_1838_0;
          st_2 <= `S_2_1201;
        end
        `S_2_1201: begin
          r4_Ch_6_870 <= insn_o_2_1840_0;
          st_2 <= `S_2_1202;
        end
        `S_2_1202: begin
          r3_Ch_3_871 <= r4_Ch_6_870;
          st_2 <= `S_2_676;
        end
        `S_2_1209: begin
          arg_192_879 <= x_15_872;
          st_2 <= `S_2_1227;
        end
        `S_2_1210: begin
          r4_e0_17_873 <= r1_ror32_2_193_883;
          st_2 <= `S_2_1212;
        end
        `S_2_1212: begin
          arg_172_884 <= x_15_872;
          st_2 <= `S_2_1240;
        end
        `S_2_1213: begin
          r6_e0_18_874 <= r1_ror32_13_173_888;
          st_2 <= `S_2_1214;
        end
        `S_2_1214: begin
          r3_e0_19_875 <= insn_o_2_1861_0;
          st_2 <= `S_2_1216;
        end
        `S_2_1216: begin
          arg_197_889 <= x_15_872;
          st_2 <= `S_2_1253;
        end
        `S_2_1217: begin
          r8_e0_20_876 <= r1_ror32_22_198_893;
          st_2 <= `S_2_1218;
        end
        `S_2_1218: begin
          r2_e0_21_877 <= insn_o_2_1869_0;
          st_2 <= `S_2_1219;
        end
        `S_2_1219: begin
          r1_e0_16_878 <= r2_e0_21_877;
          st_2 <= `S_2_693;
        end
        `S_2_1227: begin
          r3_ror32_2_194_880 <= insn_o_2_1880_0;
          st_2 <= `S_2_1230;
        end
        `S_2_1230: begin
          r6_ror32_2_195_881 <= insn_o_2_1884_0;
          st_2 <= `S_2_1231;
        end
        `S_2_1231: begin
          r2_ror32_2_196_882 <= insn_o_2_1886_0;
          st_2 <= `S_2_1232;
        end
        `S_2_1232: begin
          r1_ror32_2_193_883 <= r2_ror32_2_196_882;
          st_2 <= `S_2_1210;
        end
        `S_2_1240: begin
          r3_ror32_13_174_885 <= insn_o_2_1897_0;
          st_2 <= `S_2_1243;
        end
        `S_2_1243: begin
          r6_ror32_13_175_886 <= insn_o_2_1901_0;
          st_2 <= `S_2_1244;
        end
        `S_2_1244: begin
          r2_ror32_13_176_887 <= insn_o_2_1903_0;
          st_2 <= `S_2_1245;
        end
        `S_2_1245: begin
          r1_ror32_13_173_888 <= r2_ror32_13_176_887;
          st_2 <= `S_2_1213;
        end
        `S_2_1253: begin
          r3_ror32_22_199_890 <= insn_o_2_1914_0;
          st_2 <= `S_2_1256;
        end
        `S_2_1256: begin
          r6_ror32_22_200_891 <= insn_o_2_1918_0;
          st_2 <= `S_2_1257;
        end
        `S_2_1257: begin
          r2_ror32_22_201_892 <= insn_o_2_1920_0;
          st_2 <= `S_2_1258;
        end
        `S_2_1258: begin
          r1_ror32_22_198_893 <= r2_ror32_22_201_892;
          st_2 <= `S_2_1217;
        end
        `S_2_1264: begin
          r5_Maj_11_896 <= insn_o_2_1929_0;
          st_2 <= `S_2_1265;
        end
        `S_2_1265: begin
          r7_Maj_12_897 <= insn_o_2_1931_0;
          st_2 <= `S_2_1266;
        end
        `S_2_1266: begin
          r6_Maj_13_899 <= insn_o_2_1933_0;
          st_2 <= `S_2_1267;
        end
        `S_2_1267: begin
          r4_Maj_14_900 <= insn_o_2_1935_0;
          st_2 <= `S_2_1268;
        end
        `S_2_1268: begin
          r3_Maj_10_901 <= r4_Maj_14_900;
          st_2 <= `S_2_696;
        end
        `S_2_1275: begin
          arg_207_909 <= x_22_902;
          st_2 <= `S_2_1293;
        end
        `S_2_1276: begin
          r4_e1_24_903 <= r1_ror32_6_208_913;
          st_2 <= `S_2_1278;
        end
        `S_2_1278: begin
          arg_167_914 <= x_22_902;
          st_2 <= `S_2_1306;
        end
        `S_2_1279: begin
          r6_e1_25_904 <= r1_ror32_11_168_918;
          st_2 <= `S_2_1280;
        end
        `S_2_1280: begin
          r3_e1_26_905 <= insn_o_2_1956_0;
          st_2 <= `S_2_1282;
        end
        `S_2_1282: begin
          arg_202_919 <= x_22_902;
          st_2 <= `S_2_1319;
        end
        `S_2_1283: begin
          r8_e1_27_906 <= r1_ror32_25_203_923;
          st_2 <= `S_2_1284;
        end
        `S_2_1284: begin
          r2_e1_28_907 <= insn_o_2_1964_0;
          st_2 <= `S_2_1285;
        end
        `S_2_1285: begin
          r1_e1_23_908 <= r2_e1_28_907;
          st_2 <= `S_2_705;
        end
        `S_2_1293: begin
          r3_ror32_6_209_910 <= insn_o_2_1975_0;
          st_2 <= `S_2_1296;
        end
        `S_2_1296: begin
          r6_ror32_6_210_911 <= insn_o_2_1979_0;
          st_2 <= `S_2_1297;
        end
        `S_2_1297: begin
          r2_ror32_6_211_912 <= insn_o_2_1981_0;
          st_2 <= `S_2_1298;
        end
        `S_2_1298: begin
          r1_ror32_6_208_913 <= r2_ror32_6_211_912;
          st_2 <= `S_2_1276;
        end
        `S_2_1306: begin
          r3_ror32_11_169_915 <= insn_o_2_1992_0;
          st_2 <= `S_2_1309;
        end
        `S_2_1309: begin
          r6_ror32_11_170_916 <= insn_o_2_1996_0;
          st_2 <= `S_2_1310;
        end
        `S_2_1310: begin
          r2_ror32_11_171_917 <= insn_o_2_1998_0;
          st_2 <= `S_2_1311;
        end
        `S_2_1311: begin
          r1_ror32_11_168_918 <= r2_ror32_11_171_917;
          st_2 <= `S_2_1279;
        end
        `S_2_1319: begin
          r3_ror32_25_204_920 <= insn_o_2_2009_0;
          st_2 <= `S_2_1322;
        end
        `S_2_1322: begin
          r6_ror32_25_205_921 <= insn_o_2_2013_0;
          st_2 <= `S_2_1323;
        end
        `S_2_1323: begin
          r2_ror32_25_206_922 <= insn_o_2_2015_0;
          st_2 <= `S_2_1324;
        end
        `S_2_1324: begin
          r1_ror32_25_203_923 <= r2_ror32_25_206_922;
          st_2 <= `S_2_1283;
        end
        `S_2_1330: begin
          r6_Ch_4_926 <= insn_o_2_2024_0;
          st_2 <= `S_2_1331;
        end
        `S_2_1331: begin
          r5_Ch_5_928 <= insn_o_2_2026_0;
          st_2 <= `S_2_1332;
        end
        `S_2_1332: begin
          r4_Ch_6_929 <= insn_o_2_2028_0;
          st_2 <= `S_2_1333;
        end
        `S_2_1333: begin
          r3_Ch_3_930 <= r4_Ch_6_929;
          st_2 <= `S_2_709;
        end
        `S_2_1340: begin
          arg_192_938 <= x_15_931;
          st_2 <= `S_2_1358;
        end
        `S_2_1341: begin
          r4_e0_17_932 <= r1_ror32_2_193_942;
          st_2 <= `S_2_1343;
        end
        `S_2_1343: begin
          arg_172_943 <= x_15_931;
          st_2 <= `S_2_1371;
        end
        `S_2_1344: begin
          r6_e0_18_933 <= r1_ror32_13_173_947;
          st_2 <= `S_2_1345;
        end
        `S_2_1345: begin
          r3_e0_19_934 <= insn_o_2_2049_0;
          st_2 <= `S_2_1347;
        end
        `S_2_1347: begin
          arg_197_948 <= x_15_931;
          st_2 <= `S_2_1384;
        end
        `S_2_1348: begin
          r8_e0_20_935 <= r1_ror32_22_198_952;
          st_2 <= `S_2_1349;
        end
        `S_2_1349: begin
          r2_e0_21_936 <= insn_o_2_2057_0;
          st_2 <= `S_2_1350;
        end
        `S_2_1350: begin
          r1_e0_16_937 <= r2_e0_21_936;
          st_2 <= `S_2_726;
        end
        `S_2_1358: begin
          r3_ror32_2_194_939 <= insn_o_2_2068_0;
          st_2 <= `S_2_1361;
        end
        `S_2_1361: begin
          r6_ror32_2_195_940 <= insn_o_2_2072_0;
          st_2 <= `S_2_1362;
        end
        `S_2_1362: begin
          r2_ror32_2_196_941 <= insn_o_2_2074_0;
          st_2 <= `S_2_1363;
        end
        `S_2_1363: begin
          r1_ror32_2_193_942 <= r2_ror32_2_196_941;
          st_2 <= `S_2_1341;
        end
        `S_2_1371: begin
          r3_ror32_13_174_944 <= insn_o_2_2085_0;
          st_2 <= `S_2_1374;
        end
        `S_2_1374: begin
          r6_ror32_13_175_945 <= insn_o_2_2089_0;
          st_2 <= `S_2_1375;
        end
        `S_2_1375: begin
          r2_ror32_13_176_946 <= insn_o_2_2091_0;
          st_2 <= `S_2_1376;
        end
        `S_2_1376: begin
          r1_ror32_13_173_947 <= r2_ror32_13_176_946;
          st_2 <= `S_2_1344;
        end
        `S_2_1384: begin
          r3_ror32_22_199_949 <= insn_o_2_2102_0;
          st_2 <= `S_2_1387;
        end
        `S_2_1387: begin
          r6_ror32_22_200_950 <= insn_o_2_2106_0;
          st_2 <= `S_2_1388;
        end
        `S_2_1388: begin
          r2_ror32_22_201_951 <= insn_o_2_2108_0;
          st_2 <= `S_2_1389;
        end
        `S_2_1389: begin
          r1_ror32_22_198_952 <= r2_ror32_22_201_951;
          st_2 <= `S_2_1348;
        end
        `S_2_1395: begin
          r5_Maj_11_955 <= insn_o_2_2117_0;
          st_2 <= `S_2_1396;
        end
        `S_2_1396: begin
          r7_Maj_12_956 <= insn_o_2_2119_0;
          st_2 <= `S_2_1397;
        end
        `S_2_1397: begin
          r6_Maj_13_958 <= insn_o_2_2121_0;
          st_2 <= `S_2_1398;
        end
        `S_2_1398: begin
          r4_Maj_14_959 <= insn_o_2_2123_0;
          st_2 <= `S_2_1399;
        end
        `S_2_1399: begin
          r3_Maj_10_960 <= r4_Maj_14_959;
          st_2 <= `S_2_729;
        end
        `S_2_1406: begin
          arg_207_968 <= x_22_961;
          st_2 <= `S_2_1424;
        end
        `S_2_1407: begin
          r4_e1_24_962 <= r1_ror32_6_208_972;
          st_2 <= `S_2_1409;
        end
        `S_2_1409: begin
          arg_167_973 <= x_22_961;
          st_2 <= `S_2_1437;
        end
        `S_2_1410: begin
          r6_e1_25_963 <= r1_ror32_11_168_977;
          st_2 <= `S_2_1411;
        end
        `S_2_1411: begin
          r3_e1_26_964 <= insn_o_2_2144_0;
          st_2 <= `S_2_1413;
        end
        `S_2_1413: begin
          arg_202_978 <= x_22_961;
          st_2 <= `S_2_1450;
        end
        `S_2_1414: begin
          r8_e1_27_965 <= r1_ror32_25_203_982;
          st_2 <= `S_2_1415;
        end
        `S_2_1415: begin
          r2_e1_28_966 <= insn_o_2_2152_0;
          st_2 <= `S_2_1416;
        end
        `S_2_1416: begin
          r1_e1_23_967 <= r2_e1_28_966;
          st_2 <= `S_2_738;
        end
        `S_2_1424: begin
          r3_ror32_6_209_969 <= insn_o_2_2163_0;
          st_2 <= `S_2_1427;
        end
        `S_2_1427: begin
          r6_ror32_6_210_970 <= insn_o_2_2167_0;
          st_2 <= `S_2_1428;
        end
        `S_2_1428: begin
          r2_ror32_6_211_971 <= insn_o_2_2169_0;
          st_2 <= `S_2_1429;
        end
        `S_2_1429: begin
          r1_ror32_6_208_972 <= r2_ror32_6_211_971;
          st_2 <= `S_2_1407;
        end
        `S_2_1437: begin
          r3_ror32_11_169_974 <= insn_o_2_2180_0;
          st_2 <= `S_2_1440;
        end
        `S_2_1440: begin
          r6_ror32_11_170_975 <= insn_o_2_2184_0;
          st_2 <= `S_2_1441;
        end
        `S_2_1441: begin
          r2_ror32_11_171_976 <= insn_o_2_2186_0;
          st_2 <= `S_2_1442;
        end
        `S_2_1442: begin
          r1_ror32_11_168_977 <= r2_ror32_11_171_976;
          st_2 <= `S_2_1410;
        end
        `S_2_1450: begin
          r3_ror32_25_204_979 <= insn_o_2_2197_0;
          st_2 <= `S_2_1453;
        end
        `S_2_1453: begin
          r6_ror32_25_205_980 <= insn_o_2_2201_0;
          st_2 <= `S_2_1454;
        end
        `S_2_1454: begin
          r2_ror32_25_206_981 <= insn_o_2_2203_0;
          st_2 <= `S_2_1455;
        end
        `S_2_1455: begin
          r1_ror32_25_203_982 <= r2_ror32_25_206_981;
          st_2 <= `S_2_1414;
        end
        `S_2_1461: begin
          r6_Ch_4_985 <= insn_o_2_2212_0;
          st_2 <= `S_2_1462;
        end
        `S_2_1462: begin
          r5_Ch_5_987 <= insn_o_2_2214_0;
          st_2 <= `S_2_1463;
        end
        `S_2_1463: begin
          r4_Ch_6_988 <= insn_o_2_2216_0;
          st_2 <= `S_2_1464;
        end
        `S_2_1464: begin
          r3_Ch_3_989 <= r4_Ch_6_988;
          st_2 <= `S_2_742;
        end
        `S_2_1471: begin
          arg_192_997 <= x_15_990;
          st_2 <= `S_2_1489;
        end
        `S_2_1472: begin
          r4_e0_17_991 <= r1_ror32_2_193_1001;
          st_2 <= `S_2_1474;
        end
        `S_2_1474: begin
          arg_172_1002 <= x_15_990;
          st_2 <= `S_2_1502;
        end
        `S_2_1475: begin
          r6_e0_18_992 <= r1_ror32_13_173_1006;
          st_2 <= `S_2_1476;
        end
        `S_2_1476: begin
          r3_e0_19_993 <= insn_o_2_2237_0;
          st_2 <= `S_2_1478;
        end
        `S_2_1478: begin
          arg_197_1007 <= x_15_990;
          st_2 <= `S_2_1515;
        end
        `S_2_1479: begin
          r8_e0_20_994 <= r1_ror32_22_198_1011;
          st_2 <= `S_2_1480;
        end
        `S_2_1480: begin
          r2_e0_21_995 <= insn_o_2_2245_0;
          st_2 <= `S_2_1481;
        end
        `S_2_1481: begin
          r1_e0_16_996 <= r2_e0_21_995;
          st_2 <= `S_2_759;
        end
        `S_2_1489: begin
          r3_ror32_2_194_998 <= insn_o_2_2256_0;
          st_2 <= `S_2_1492;
        end
        `S_2_1492: begin
          r6_ror32_2_195_999 <= insn_o_2_2260_0;
          st_2 <= `S_2_1493;
        end
        `S_2_1493: begin
          r2_ror32_2_196_1000 <= insn_o_2_2262_0;
          st_2 <= `S_2_1494;
        end
        `S_2_1494: begin
          r1_ror32_2_193_1001 <= r2_ror32_2_196_1000;
          st_2 <= `S_2_1472;
        end
        `S_2_1502: begin
          r3_ror32_13_174_1003 <= insn_o_2_2273_0;
          st_2 <= `S_2_1505;
        end
        `S_2_1505: begin
          r6_ror32_13_175_1004 <= insn_o_2_2277_0;
          st_2 <= `S_2_1506;
        end
        `S_2_1506: begin
          r2_ror32_13_176_1005 <= insn_o_2_2279_0;
          st_2 <= `S_2_1507;
        end
        `S_2_1507: begin
          r1_ror32_13_173_1006 <= r2_ror32_13_176_1005;
          st_2 <= `S_2_1475;
        end
        `S_2_1515: begin
          r3_ror32_22_199_1008 <= insn_o_2_2290_0;
          st_2 <= `S_2_1518;
        end
        `S_2_1518: begin
          r6_ror32_22_200_1009 <= insn_o_2_2294_0;
          st_2 <= `S_2_1519;
        end
        `S_2_1519: begin
          r2_ror32_22_201_1010 <= insn_o_2_2296_0;
          st_2 <= `S_2_1520;
        end
        `S_2_1520: begin
          r1_ror32_22_198_1011 <= r2_ror32_22_201_1010;
          st_2 <= `S_2_1479;
        end
        `S_2_1526: begin
          r5_Maj_11_1014 <= insn_o_2_2305_0;
          st_2 <= `S_2_1527;
        end
        `S_2_1527: begin
          r7_Maj_12_1015 <= insn_o_2_2307_0;
          st_2 <= `S_2_1528;
        end
        `S_2_1528: begin
          r6_Maj_13_1017 <= insn_o_2_2309_0;
          st_2 <= `S_2_1529;
        end
        `S_2_1529: begin
          r4_Maj_14_1018 <= insn_o_2_2311_0;
          st_2 <= `S_2_1530;
        end
        `S_2_1530: begin
          r3_Maj_10_1019 <= r4_Maj_14_1018;
          st_2 <= `S_2_762;
        end
        `S_2_1537: begin
          arg_207_1027 <= x_22_1020;
          st_2 <= `S_2_1555;
        end
        `S_2_1538: begin
          r4_e1_24_1021 <= r1_ror32_6_208_1031;
          st_2 <= `S_2_1540;
        end
        `S_2_1540: begin
          arg_167_1032 <= x_22_1020;
          st_2 <= `S_2_1568;
        end
        `S_2_1541: begin
          r6_e1_25_1022 <= r1_ror32_11_168_1036;
          st_2 <= `S_2_1542;
        end
        `S_2_1542: begin
          r3_e1_26_1023 <= insn_o_2_2332_0;
          st_2 <= `S_2_1544;
        end
        `S_2_1544: begin
          arg_202_1037 <= x_22_1020;
          st_2 <= `S_2_1581;
        end
        `S_2_1545: begin
          r8_e1_27_1024 <= r1_ror32_25_203_1041;
          st_2 <= `S_2_1546;
        end
        `S_2_1546: begin
          r2_e1_28_1025 <= insn_o_2_2340_0;
          st_2 <= `S_2_1547;
        end
        `S_2_1547: begin
          r1_e1_23_1026 <= r2_e1_28_1025;
          st_2 <= `S_2_771;
        end
        `S_2_1555: begin
          r3_ror32_6_209_1028 <= insn_o_2_2351_0;
          st_2 <= `S_2_1558;
        end
        `S_2_1558: begin
          r6_ror32_6_210_1029 <= insn_o_2_2355_0;
          st_2 <= `S_2_1559;
        end
        `S_2_1559: begin
          r2_ror32_6_211_1030 <= insn_o_2_2357_0;
          st_2 <= `S_2_1560;
        end
        `S_2_1560: begin
          r1_ror32_6_208_1031 <= r2_ror32_6_211_1030;
          st_2 <= `S_2_1538;
        end
        `S_2_1568: begin
          r3_ror32_11_169_1033 <= insn_o_2_2368_0;
          st_2 <= `S_2_1571;
        end
        `S_2_1571: begin
          r6_ror32_11_170_1034 <= insn_o_2_2372_0;
          st_2 <= `S_2_1572;
        end
        `S_2_1572: begin
          r2_ror32_11_171_1035 <= insn_o_2_2374_0;
          st_2 <= `S_2_1573;
        end
        `S_2_1573: begin
          r1_ror32_11_168_1036 <= r2_ror32_11_171_1035;
          st_2 <= `S_2_1541;
        end
        `S_2_1581: begin
          r3_ror32_25_204_1038 <= insn_o_2_2385_0;
          st_2 <= `S_2_1584;
        end
        `S_2_1584: begin
          r6_ror32_25_205_1039 <= insn_o_2_2389_0;
          st_2 <= `S_2_1585;
        end
        `S_2_1585: begin
          r2_ror32_25_206_1040 <= insn_o_2_2391_0;
          st_2 <= `S_2_1586;
        end
        `S_2_1586: begin
          r1_ror32_25_203_1041 <= r2_ror32_25_206_1040;
          st_2 <= `S_2_1545;
        end
        `S_2_1592: begin
          r6_Ch_4_1044 <= insn_o_2_2400_0;
          st_2 <= `S_2_1593;
        end
        `S_2_1593: begin
          r5_Ch_5_1046 <= insn_o_2_2402_0;
          st_2 <= `S_2_1594;
        end
        `S_2_1594: begin
          r4_Ch_6_1047 <= insn_o_2_2404_0;
          st_2 <= `S_2_1595;
        end
        `S_2_1595: begin
          r3_Ch_3_1048 <= r4_Ch_6_1047;
          st_2 <= `S_2_775;
        end
        `S_2_1602: begin
          arg_192_1056 <= x_15_1049;
          st_2 <= `S_2_1620;
        end
        `S_2_1603: begin
          r4_e0_17_1050 <= r1_ror32_2_193_1060;
          st_2 <= `S_2_1605;
        end
        `S_2_1605: begin
          arg_172_1061 <= x_15_1049;
          st_2 <= `S_2_1633;
        end
        `S_2_1606: begin
          r6_e0_18_1051 <= r1_ror32_13_173_1065;
          st_2 <= `S_2_1607;
        end
        `S_2_1607: begin
          r3_e0_19_1052 <= insn_o_2_2425_0;
          st_2 <= `S_2_1609;
        end
        `S_2_1609: begin
          arg_197_1066 <= x_15_1049;
          st_2 <= `S_2_1646;
        end
        `S_2_1610: begin
          r8_e0_20_1053 <= r1_ror32_22_198_1070;
          st_2 <= `S_2_1611;
        end
        `S_2_1611: begin
          r2_e0_21_1054 <= insn_o_2_2433_0;
          st_2 <= `S_2_1612;
        end
        `S_2_1612: begin
          r1_e0_16_1055 <= r2_e0_21_1054;
          st_2 <= `S_2_792;
        end
        `S_2_1620: begin
          r3_ror32_2_194_1057 <= insn_o_2_2444_0;
          st_2 <= `S_2_1623;
        end
        `S_2_1623: begin
          r6_ror32_2_195_1058 <= insn_o_2_2448_0;
          st_2 <= `S_2_1624;
        end
        `S_2_1624: begin
          r2_ror32_2_196_1059 <= insn_o_2_2450_0;
          st_2 <= `S_2_1625;
        end
        `S_2_1625: begin
          r1_ror32_2_193_1060 <= r2_ror32_2_196_1059;
          st_2 <= `S_2_1603;
        end
        `S_2_1633: begin
          r3_ror32_13_174_1062 <= insn_o_2_2461_0;
          st_2 <= `S_2_1636;
        end
        `S_2_1636: begin
          r6_ror32_13_175_1063 <= insn_o_2_2465_0;
          st_2 <= `S_2_1637;
        end
        `S_2_1637: begin
          r2_ror32_13_176_1064 <= insn_o_2_2467_0;
          st_2 <= `S_2_1638;
        end
        `S_2_1638: begin
          r1_ror32_13_173_1065 <= r2_ror32_13_176_1064;
          st_2 <= `S_2_1606;
        end
        `S_2_1646: begin
          r3_ror32_22_199_1067 <= insn_o_2_2478_0;
          st_2 <= `S_2_1649;
        end
        `S_2_1649: begin
          r6_ror32_22_200_1068 <= insn_o_2_2482_0;
          st_2 <= `S_2_1650;
        end
        `S_2_1650: begin
          r2_ror32_22_201_1069 <= insn_o_2_2484_0;
          st_2 <= `S_2_1651;
        end
        `S_2_1651: begin
          r1_ror32_22_198_1070 <= r2_ror32_22_201_1069;
          st_2 <= `S_2_1610;
        end
        `S_2_1657: begin
          r5_Maj_11_1073 <= insn_o_2_2493_0;
          st_2 <= `S_2_1658;
        end
        `S_2_1658: begin
          r7_Maj_12_1074 <= insn_o_2_2495_0;
          st_2 <= `S_2_1659;
        end
        `S_2_1659: begin
          r6_Maj_13_1076 <= insn_o_2_2497_0;
          st_2 <= `S_2_1660;
        end
        `S_2_1660: begin
          r4_Maj_14_1077 <= insn_o_2_2499_0;
          st_2 <= `S_2_1661;
        end
        `S_2_1661: begin
          r3_Maj_10_1078 <= r4_Maj_14_1077;
          st_2 <= `S_2_795;
        end
        `S_2_1668: begin
          arg_207_1086 <= x_22_1079;
          st_2 <= `S_2_1686;
        end
        `S_2_1669: begin
          r4_e1_24_1080 <= r1_ror32_6_208_1090;
          st_2 <= `S_2_1671;
        end
        `S_2_1671: begin
          arg_167_1091 <= x_22_1079;
          st_2 <= `S_2_1699;
        end
        `S_2_1672: begin
          r6_e1_25_1081 <= r1_ror32_11_168_1095;
          st_2 <= `S_2_1673;
        end
        `S_2_1673: begin
          r3_e1_26_1082 <= insn_o_2_2520_0;
          st_2 <= `S_2_1675;
        end
        `S_2_1675: begin
          arg_202_1096 <= x_22_1079;
          st_2 <= `S_2_1712;
        end
        `S_2_1676: begin
          r8_e1_27_1083 <= r1_ror32_25_203_1100;
          st_2 <= `S_2_1677;
        end
        `S_2_1677: begin
          r2_e1_28_1084 <= insn_o_2_2528_0;
          st_2 <= `S_2_1678;
        end
        `S_2_1678: begin
          r1_e1_23_1085 <= r2_e1_28_1084;
          st_2 <= `S_2_804;
        end
        `S_2_1686: begin
          r3_ror32_6_209_1087 <= insn_o_2_2539_0;
          st_2 <= `S_2_1689;
        end
        `S_2_1689: begin
          r6_ror32_6_210_1088 <= insn_o_2_2543_0;
          st_2 <= `S_2_1690;
        end
        `S_2_1690: begin
          r2_ror32_6_211_1089 <= insn_o_2_2545_0;
          st_2 <= `S_2_1691;
        end
        `S_2_1691: begin
          r1_ror32_6_208_1090 <= r2_ror32_6_211_1089;
          st_2 <= `S_2_1669;
        end
        `S_2_1699: begin
          r3_ror32_11_169_1092 <= insn_o_2_2556_0;
          st_2 <= `S_2_1702;
        end
        `S_2_1702: begin
          r6_ror32_11_170_1093 <= insn_o_2_2560_0;
          st_2 <= `S_2_1703;
        end
        `S_2_1703: begin
          r2_ror32_11_171_1094 <= insn_o_2_2562_0;
          st_2 <= `S_2_1704;
        end
        `S_2_1704: begin
          r1_ror32_11_168_1095 <= r2_ror32_11_171_1094;
          st_2 <= `S_2_1672;
        end
        `S_2_1712: begin
          r3_ror32_25_204_1097 <= insn_o_2_2573_0;
          st_2 <= `S_2_1715;
        end
        `S_2_1715: begin
          r6_ror32_25_205_1098 <= insn_o_2_2577_0;
          st_2 <= `S_2_1716;
        end
        `S_2_1716: begin
          r2_ror32_25_206_1099 <= insn_o_2_2579_0;
          st_2 <= `S_2_1717;
        end
        `S_2_1717: begin
          r1_ror32_25_203_1100 <= r2_ror32_25_206_1099;
          st_2 <= `S_2_1676;
        end
        `S_2_1723: begin
          r6_Ch_4_1103 <= insn_o_2_2588_0;
          st_2 <= `S_2_1724;
        end
        `S_2_1724: begin
          r5_Ch_5_1105 <= insn_o_2_2590_0;
          st_2 <= `S_2_1725;
        end
        `S_2_1725: begin
          r4_Ch_6_1106 <= insn_o_2_2592_0;
          st_2 <= `S_2_1726;
        end
        `S_2_1726: begin
          r3_Ch_3_1107 <= r4_Ch_6_1106;
          st_2 <= `S_2_808;
        end
        `S_2_1733: begin
          arg_192_1115 <= x_15_1108;
          st_2 <= `S_2_1751;
        end
        `S_2_1734: begin
          r4_e0_17_1109 <= r1_ror32_2_193_1119;
          st_2 <= `S_2_1736;
        end
        `S_2_1736: begin
          arg_172_1120 <= x_15_1108;
          st_2 <= `S_2_1764;
        end
        `S_2_1737: begin
          r6_e0_18_1110 <= r1_ror32_13_173_1124;
          st_2 <= `S_2_1738;
        end
        `S_2_1738: begin
          r3_e0_19_1111 <= insn_o_2_2613_0;
          st_2 <= `S_2_1740;
        end
        `S_2_1740: begin
          arg_197_1125 <= x_15_1108;
          st_2 <= `S_2_1777;
        end
        `S_2_1741: begin
          r8_e0_20_1112 <= r1_ror32_22_198_1129;
          st_2 <= `S_2_1742;
        end
        `S_2_1742: begin
          r2_e0_21_1113 <= insn_o_2_2621_0;
          st_2 <= `S_2_1743;
        end
        `S_2_1743: begin
          r1_e0_16_1114 <= r2_e0_21_1113;
          st_2 <= `S_2_825;
        end
        `S_2_1751: begin
          r3_ror32_2_194_1116 <= insn_o_2_2632_0;
          st_2 <= `S_2_1754;
        end
        `S_2_1754: begin
          r6_ror32_2_195_1117 <= insn_o_2_2636_0;
          st_2 <= `S_2_1755;
        end
        `S_2_1755: begin
          r2_ror32_2_196_1118 <= insn_o_2_2638_0;
          st_2 <= `S_2_1756;
        end
        `S_2_1756: begin
          r1_ror32_2_193_1119 <= r2_ror32_2_196_1118;
          st_2 <= `S_2_1734;
        end
        `S_2_1764: begin
          r3_ror32_13_174_1121 <= insn_o_2_2649_0;
          st_2 <= `S_2_1767;
        end
        `S_2_1767: begin
          r6_ror32_13_175_1122 <= insn_o_2_2653_0;
          st_2 <= `S_2_1768;
        end
        `S_2_1768: begin
          r2_ror32_13_176_1123 <= insn_o_2_2655_0;
          st_2 <= `S_2_1769;
        end
        `S_2_1769: begin
          r1_ror32_13_173_1124 <= r2_ror32_13_176_1123;
          st_2 <= `S_2_1737;
        end
        `S_2_1777: begin
          r3_ror32_22_199_1126 <= insn_o_2_2666_0;
          st_2 <= `S_2_1780;
        end
        `S_2_1780: begin
          r6_ror32_22_200_1127 <= insn_o_2_2670_0;
          st_2 <= `S_2_1781;
        end
        `S_2_1781: begin
          r2_ror32_22_201_1128 <= insn_o_2_2672_0;
          st_2 <= `S_2_1782;
        end
        `S_2_1782: begin
          r1_ror32_22_198_1129 <= r2_ror32_22_201_1128;
          st_2 <= `S_2_1741;
        end
        `S_2_1788: begin
          r5_Maj_11_1132 <= insn_o_2_2681_0;
          st_2 <= `S_2_1789;
        end
        `S_2_1789: begin
          r7_Maj_12_1133 <= insn_o_2_2683_0;
          st_2 <= `S_2_1790;
        end
        `S_2_1790: begin
          r6_Maj_13_1135 <= insn_o_2_2685_0;
          st_2 <= `S_2_1791;
        end
        `S_2_1791: begin
          r4_Maj_14_1136 <= insn_o_2_2687_0;
          st_2 <= `S_2_1792;
        end
        `S_2_1792: begin
          r3_Maj_10_1137 <= r4_Maj_14_1136;
          st_2 <= `S_2_828;
        end
        `S_2_1799: begin
          arg_207_1145 <= x_22_1138;
          st_2 <= `S_2_1817;
        end
        `S_2_1800: begin
          r4_e1_24_1139 <= r1_ror32_6_208_1149;
          st_2 <= `S_2_1802;
        end
        `S_2_1802: begin
          arg_167_1150 <= x_22_1138;
          st_2 <= `S_2_1830;
        end
        `S_2_1803: begin
          r6_e1_25_1140 <= r1_ror32_11_168_1154;
          st_2 <= `S_2_1804;
        end
        `S_2_1804: begin
          r3_e1_26_1141 <= insn_o_2_2708_0;
          st_2 <= `S_2_1806;
        end
        `S_2_1806: begin
          arg_202_1155 <= x_22_1138;
          st_2 <= `S_2_1843;
        end
        `S_2_1807: begin
          r8_e1_27_1142 <= r1_ror32_25_203_1159;
          st_2 <= `S_2_1808;
        end
        `S_2_1808: begin
          r2_e1_28_1143 <= insn_o_2_2716_0;
          st_2 <= `S_2_1809;
        end
        `S_2_1809: begin
          r1_e1_23_1144 <= r2_e1_28_1143;
          st_2 <= `S_2_837;
        end
        `S_2_1817: begin
          r3_ror32_6_209_1146 <= insn_o_2_2727_0;
          st_2 <= `S_2_1820;
        end
        `S_2_1820: begin
          r6_ror32_6_210_1147 <= insn_o_2_2731_0;
          st_2 <= `S_2_1821;
        end
        `S_2_1821: begin
          r2_ror32_6_211_1148 <= insn_o_2_2733_0;
          st_2 <= `S_2_1822;
        end
        `S_2_1822: begin
          r1_ror32_6_208_1149 <= r2_ror32_6_211_1148;
          st_2 <= `S_2_1800;
        end
        `S_2_1830: begin
          r3_ror32_11_169_1151 <= insn_o_2_2744_0;
          st_2 <= `S_2_1833;
        end
        `S_2_1833: begin
          r6_ror32_11_170_1152 <= insn_o_2_2748_0;
          st_2 <= `S_2_1834;
        end
        `S_2_1834: begin
          r2_ror32_11_171_1153 <= insn_o_2_2750_0;
          st_2 <= `S_2_1835;
        end
        `S_2_1835: begin
          r1_ror32_11_168_1154 <= r2_ror32_11_171_1153;
          st_2 <= `S_2_1803;
        end
        `S_2_1843: begin
          r3_ror32_25_204_1156 <= insn_o_2_2761_0;
          st_2 <= `S_2_1846;
        end
        `S_2_1846: begin
          r6_ror32_25_205_1157 <= insn_o_2_2765_0;
          st_2 <= `S_2_1847;
        end
        `S_2_1847: begin
          r2_ror32_25_206_1158 <= insn_o_2_2767_0;
          st_2 <= `S_2_1848;
        end
        `S_2_1848: begin
          r1_ror32_25_203_1159 <= r2_ror32_25_206_1158;
          st_2 <= `S_2_1807;
        end
        `S_2_1854: begin
          r6_Ch_4_1162 <= insn_o_2_2776_0;
          st_2 <= `S_2_1855;
        end
        `S_2_1855: begin
          r5_Ch_5_1164 <= insn_o_2_2778_0;
          st_2 <= `S_2_1856;
        end
        `S_2_1856: begin
          r4_Ch_6_1165 <= insn_o_2_2780_0;
          st_2 <= `S_2_1857;
        end
        `S_2_1857: begin
          r3_Ch_3_1166 <= r4_Ch_6_1165;
          st_2 <= `S_2_841;
        end
        `S_2_1864: begin
          arg_192_1174 <= x_15_1167;
          st_2 <= `S_2_1882;
        end
        `S_2_1865: begin
          r4_e0_17_1168 <= r1_ror32_2_193_1178;
          st_2 <= `S_2_1867;
        end
        `S_2_1867: begin
          arg_172_1179 <= x_15_1167;
          st_2 <= `S_2_1895;
        end
        `S_2_1868: begin
          r6_e0_18_1169 <= r1_ror32_13_173_1183;
          st_2 <= `S_2_1869;
        end
        `S_2_1869: begin
          r3_e0_19_1170 <= insn_o_2_2801_0;
          st_2 <= `S_2_1871;
        end
        `S_2_1871: begin
          arg_197_1184 <= x_15_1167;
          st_2 <= `S_2_1908;
        end
        `S_2_1872: begin
          r8_e0_20_1171 <= r1_ror32_22_198_1188;
          st_2 <= `S_2_1873;
        end
        `S_2_1873: begin
          r2_e0_21_1172 <= insn_o_2_2809_0;
          st_2 <= `S_2_1874;
        end
        `S_2_1874: begin
          r1_e0_16_1173 <= r2_e0_21_1172;
          st_2 <= `S_2_858;
        end
        `S_2_1882: begin
          r3_ror32_2_194_1175 <= insn_o_2_2820_0;
          st_2 <= `S_2_1885;
        end
        `S_2_1885: begin
          r6_ror32_2_195_1176 <= insn_o_2_2824_0;
          st_2 <= `S_2_1886;
        end
        `S_2_1886: begin
          r2_ror32_2_196_1177 <= insn_o_2_2826_0;
          st_2 <= `S_2_1887;
        end
        `S_2_1887: begin
          r1_ror32_2_193_1178 <= r2_ror32_2_196_1177;
          st_2 <= `S_2_1865;
        end
        `S_2_1895: begin
          r3_ror32_13_174_1180 <= insn_o_2_2837_0;
          st_2 <= `S_2_1898;
        end
        `S_2_1898: begin
          r6_ror32_13_175_1181 <= insn_o_2_2841_0;
          st_2 <= `S_2_1899;
        end
        `S_2_1899: begin
          r2_ror32_13_176_1182 <= insn_o_2_2843_0;
          st_2 <= `S_2_1900;
        end
        `S_2_1900: begin
          r1_ror32_13_173_1183 <= r2_ror32_13_176_1182;
          st_2 <= `S_2_1868;
        end
        `S_2_1908: begin
          r3_ror32_22_199_1185 <= insn_o_2_2854_0;
          st_2 <= `S_2_1911;
        end
        `S_2_1911: begin
          r6_ror32_22_200_1186 <= insn_o_2_2858_0;
          st_2 <= `S_2_1912;
        end
        `S_2_1912: begin
          r2_ror32_22_201_1187 <= insn_o_2_2860_0;
          st_2 <= `S_2_1913;
        end
        `S_2_1913: begin
          r1_ror32_22_198_1188 <= r2_ror32_22_201_1187;
          st_2 <= `S_2_1872;
        end
        `S_2_1919: begin
          r5_Maj_11_1191 <= insn_o_2_2869_0;
          st_2 <= `S_2_1920;
        end
        `S_2_1920: begin
          r7_Maj_12_1192 <= insn_o_2_2871_0;
          st_2 <= `S_2_1921;
        end
        `S_2_1921: begin
          r6_Maj_13_1194 <= insn_o_2_2873_0;
          st_2 <= `S_2_1922;
        end
        `S_2_1922: begin
          r4_Maj_14_1195 <= insn_o_2_2875_0;
          st_2 <= `S_2_1923;
        end
        `S_2_1923: begin
          r3_Maj_10_1196 <= r4_Maj_14_1195;
          st_2 <= `S_2_861;
        end
      endcase
    end
  end
  SRAM_4_32_2 SRAM_4_32_2_inst_2_125(.clk(clk), .rst(rst), .addr_0_i(mem_1_2_125_p0_addr), .rdata_0_o(mem_1_2_125_p0_rdata), .wdata_0_i(mem_1_2_125_p0_wdata), .write_en_0_i(mem_1_2_125_p0_wen), .addr_1_i(mem_1_2_125_p1_addr), .rdata_1_o(mem_1_2_125_p1_rdata), .wdata_1_i(mem_1_2_125_p1_wdata), .write_en_1_i(mem_1_2_125_p1_wen));
  axi_master_controller_a4rd32 inst_2_126_axi_master_controller_a4rd32(.clk(clk), .rst(rst), .sram_addr(mem_1_2_125_p1_addr), .sram_wdata(mem_1_2_125_p1_wdata), .sram_rdata(mem_1_2_125_p1_rdata), .sram_wen(mem_1_2_125_p1_wen), .sram_EXCLUSIVE(1), .sram_req(/*not connected*/), .sram_ack(1), .addr(axi_addr2_126), .wen(axi_wen2_126), .req(axi_req2_126), .len(axi_len2_126), .start(axi_start2_126), .ack(axi_ack2_126) , .ARADDR(buf_ARADDR), .ARVALID(buf_ARVALID), .ARREADY(buf_ARREADY), .ARLEN(buf_ARLEN), .ARSIZE(buf_ARSIZE), .RVALID(buf_RVALID), .RDATA(buf_RDATA), .RREADY(buf_RREADY), .RLAST(buf_RLAST), .AWADDR(buf_AWADDR), .AWVALID(buf_AWVALID), .AWREADY(buf_AWREADY), .AWLEN(buf_AWLEN), .AWSIZE(buf_AWSIZE), .WVALID(buf_WVALID), .WREADY(buf_WREADY), .WDATA(buf_WDATA), .WLAST(buf_WLAST), .BVALID(buf_BVALID), .BREADY(buf_BREADY), .BRESP(buf_BRESP));
  SRAM_3_32 SRAM_3_32_inst_2(.clk(clk), .rst(rst), .addr_i(sram_addr_2), .rdata_o(sram_rdata_2), .wdata_i(sram_wdata_2), .write_en_i(sram_wdata_en_2));
  SRAM_6_32 SRAM_6_32_inst_222(.clk(clk), .rst(rst), .addr_i(sram_addr_222), .rdata_o(sram_rdata_222), .wdata_i(sram_wdata_222), .write_en_i(sram_wdata_en_222));
  SRAM_6_32 SRAM_6_32_inst_223(.clk(clk), .rst(rst), .addr_i(sram_addr_223), .rdata_o(sram_rdata_223), .wdata_i(sram_wdata_223), .write_en_i(sram_wdata_en_223));

endmodule // main
module sha256(clk, rst, buf_ARADDR, buf_ARVALID, buf_ARREADY, buf_ARLEN, buf_ARSIZE, buf_RVALID, buf_RDATA, buf_RREADY, buf_RLAST, buf_AWADDR, buf_AWVALID, buf_AWREADY, buf_AWLEN, buf_AWSIZE, buf_WVALID, buf_WREADY, buf_WDATA, buf_WLAST, buf_BVALID, buf_BREADY, buf_BRESP, sha256_req_valid, sha256_req_ready, sha256_req_busy, sha256_res_valid, sha256_res_ready, sha256_req_0, sha256_req_1, sha256_res_0);
  input clk;
  input rst;
  output [31:0] buf_ARADDR;
  output buf_ARVALID;
  input buf_ARREADY;
  output [7:0] buf_ARLEN;
  output [2:0] buf_ARSIZE;
  input buf_RVALID;
  input [31:0] buf_RDATA;
  output buf_RREADY;
  input buf_RLAST;
  output [31:0] buf_AWADDR;
  output buf_AWVALID;
  input buf_AWREADY;
  output [7:0] buf_AWLEN;
  output [2:0] buf_AWSIZE;
  output buf_WVALID;
  input buf_WREADY;
  output [31:0] buf_WDATA;
  output buf_WLAST;
  input buf_BVALID;
  output buf_BREADY;
  input [1:0] buf_BRESP;
  input sha256_req_valid;
  output sha256_req_ready;
  output sha256_req_busy;
  output sha256_res_valid;
  input sha256_res_ready;
  input [31:0] sha256_req_0;
  input [31:0] sha256_req_1;
  output [255:0] sha256_res_0;
  main main_inst(.clk(clk), .rst(rst), .buf_ARADDR(buf_ARADDR), .buf_ARVALID(buf_ARVALID), .buf_ARREADY(buf_ARREADY), .buf_ARLEN(buf_ARLEN), .buf_ARSIZE(buf_ARSIZE), .buf_RVALID(buf_RVALID), .buf_RDATA(buf_RDATA), .buf_RREADY(buf_RREADY), .buf_RLAST(buf_RLAST), .buf_AWADDR(buf_AWADDR), .buf_AWVALID(buf_AWVALID), .buf_AWREADY(buf_AWREADY), .buf_AWLEN(buf_AWLEN), .buf_AWSIZE(buf_AWSIZE), .buf_WVALID(buf_WVALID), .buf_WREADY(buf_WREADY), .buf_WDATA(buf_WDATA), .buf_WLAST(buf_WLAST), .buf_BVALID(buf_BVALID), .buf_BREADY(buf_BREADY), .buf_BRESP(buf_BRESP), .sha256_req_valid(sha256_req_valid), .sha256_req_ready(sha256_req_ready), .sha256_req_busy(sha256_req_busy), .sha256_res_valid(sha256_res_valid), .sha256_res_ready(sha256_res_ready), .sha256_req_0(sha256_req_0), .sha256_req_1(sha256_req_1), .sha256_res_0(sha256_res_0));
endmodule
